module i2c(
    pi133,
    pi026,
    pi043,
    pi019,
    pi083,
    pi005,
    pi033,
    pi075,
    pi067,
    pi039,
    pi136,
    pi060,
    pi025,
    pi036,
    pi003,
    pi086,
    pi138,
    pi144,
    pi130,
    pi098,
    pi121,
    pi040,
    pi055,
    pi110,
    pi120,
    pi099,
    pi058,
    pi031,
    pi032,
    pi014,
    pi141,
    pi089,
    pi076,
    pi088,
    pi016,
    pi022,
    pi007,
    pi106,
    pi056,
    pi142,
    pi087,
    pi135,
    pi140,
    pi128,
    pi013,
    pi035,
    pi077,
    pi070,
    pi050,
    pi051,
    pi139,
    pi132,
    pi008,
    pi009,
    pi029,
    pi038,
    pi001,
    pi028,
    pi063,
    pi092,
    pi048,
    pi093,
    pi062,
    pi052,
    pi116,
    pi119,
    pi024,
    pi125,
    pi081,
    pi124,
    pi103,
    pi127,
    pi082,
    pi080,
    pi107,
    pi046,
    pi078,
    pi006,
    pi030,
    pi015,
    pi049,
    pi118,
    pi146,
    pi042,
    pi053,
    pi018,
    pi057,
    pi122,
    pi102,
    pi111,
    pi000,
    pi061,
    pi112,
    pi115,
    pi065,
    pi097,
    pi034,
    pi101,
    pi113,
    pi023,
    pi143,
    pi021,
    pi085,
    pi054,
    pi126,
    pi131,
    pi123,
    pi129,
    pi059,
    pi145,
    pi066,
    pi134,
    pi041,
    pi068,
    pi064,
    pi011,
    pi002,
    pi100,
    pi045,
    pi117,
    pi084,
    pi004,
    pi104,
    pi105,
    pi114,
    pi096,
    pi017,
    pi020,
    pi095,
    pi091,
    pi074,
    pi073,
    pi044,
    pi037,
    pi079,
    pi090,
    pi010,
    pi047,
    pi109,
    pi071,
    pi072,
    pi108,
    pi137,
    pi012,
    pi069,
    pi094,
    pi027,
    po120,
    po073,
    po070,
    po096,
    po066,
    po129,
    po126,
    po003,
    po040,
    po131,
    po140,
    po104,
    po127,
    po034,
    po137,
    po004,
    po117,
    po098,
    po124,
    po036,
    po084,
    po035,
    po042,
    po128,
    po043,
    po021,
    po006,
    po080,
    po101,
    po062,
    po122,
    po123,
    po057,
    po029,
    po055,
    po050,
    po069,
    po045,
    po059,
    po116,
    po054,
    po038,
    po089,
    po076,
    po068,
    po056,
    po005,
    po082,
    po135,
    po058,
    po072,
    po139,
    po086,
    po044,
    po060,
    po094,
    po078,
    po092,
    po018,
    po091,
    po010,
    po012,
    po100,
    po015,
    po099,
    po053,
    po049,
    po039,
    po108,
    po077,
    po011,
    po028,
    po002,
    po032,
    po103,
    po026,
    po130,
    po067,
    po107,
    po081,
    po020,
    po061,
    po047,
    po134,
    po008,
    po016,
    po112,
    po102,
    po074,
    po090,
    po065,
    po023,
    po111,
    po083,
    po110,
    po033,
    po030,
    po125,
    po048,
    po071,
    po017,
    po114,
    po022,
    po024,
    po079,
    po085,
    po113,
    po118,
    po075,
    po031,
    po037,
    po027,
    po138,
    po133,
    po105,
    po025,
    po141,
    po041,
    po064,
    po009,
    po013,
    po093,
    po007,
    po088,
    po000,
    po052,
    po097,
    po014,
    po087,
    po095,
    po109,
    po121,
    po046,
    po051,
    po136,
    po119,
    po001,
    po132,
    po063,
    po106,
    po115,
    po019);
    input pi133;
    input pi026;
    input pi043;
    input pi019;
    input pi083;
    input pi005;
    input pi033;
    input pi075;
    input pi067;
    input pi039;
    input pi136;
    input pi060;
    input pi025;
    input pi036;
    input pi003;
    input pi086;
    input pi138;
    input pi144;
    input pi130;
    input pi098;
    input pi121;
    input pi040;
    input pi055;
    input pi110;
    input pi120;
    input pi099;
    input pi058;
    input pi031;
    input pi032;
    input pi014;
    input pi141;
    input pi089;
    input pi076;
    input pi088;
    input pi016;
    input pi022;
    input pi007;
    input pi106;
    input pi056;
    input pi142;
    input pi087;
    input pi135;
    input pi140;
    input pi128;
    input pi013;
    input pi035;
    input pi077;
    input pi070;
    input pi050;
    input pi051;
    input pi139;
    input pi132;
    input pi008;
    input pi009;
    input pi029;
    input pi038;
    input pi001;
    input pi028;
    input pi063;
    input pi092;
    input pi048;
    input pi093;
    input pi062;
    input pi052;
    input pi116;
    input pi119;
    input pi024;
    input pi125;
    input pi081;
    input pi124;
    input pi103;
    input pi127;
    input pi082;
    input pi080;
    input pi107;
    input pi046;
    input pi078;
    input pi006;
    input pi030;
    input pi015;
    input pi049;
    input pi118;
    input pi146;
    input pi042;
    input pi053;
    input pi018;
    input pi057;
    input pi122;
    input pi102;
    input pi111;
    input pi000;
    input pi061;
    input pi112;
    input pi115;
    input pi065;
    input pi097;
    input pi034;
    input pi101;
    input pi113;
    input pi023;
    input pi143;
    input pi021;
    input pi085;
    input pi054;
    input pi126;
    input pi131;
    input pi123;
    input pi129;
    input pi059;
    input pi145;
    input pi066;
    input pi134;
    input pi041;
    input pi068;
    input pi064;
    input pi011;
    input pi002;
    input pi100;
    input pi045;
    input pi117;
    input pi084;
    input pi004;
    input pi104;
    input pi105;
    input pi114;
    input pi096;
    input pi017;
    input pi020;
    input pi095;
    input pi091;
    input pi074;
    input pi073;
    input pi044;
    input pi037;
    input pi079;
    input pi090;
    input pi010;
    input pi047;
    input pi109;
    input pi071;
    input pi072;
    input pi108;
    input pi137;
    input pi012;
    input pi069;
    input pi094;
    input pi027;
    output po120;
    output po073;
    output po070;
    output po096;
    output po066;
    output po129;
    output po126;
    output po003;
    output po040;
    output po131;
    output po140;
    output po104;
    output po127;
    output po034;
    output po137;
    output po004;
    output po117;
    output po098;
    output po124;
    output po036;
    output po084;
    output po035;
    output po042;
    output po128;
    output po043;
    output po021;
    output po006;
    output po080;
    output po101;
    output po062;
    output po122;
    output po123;
    output po057;
    output po029;
    output po055;
    output po050;
    output po069;
    output po045;
    output po059;
    output po116;
    output po054;
    output po038;
    output po089;
    output po076;
    output po068;
    output po056;
    output po005;
    output po082;
    output po135;
    output po058;
    output po072;
    output po139;
    output po086;
    output po044;
    output po060;
    output po094;
    output po078;
    output po092;
    output po018;
    output po091;
    output po010;
    output po012;
    output po100;
    output po015;
    output po099;
    output po053;
    output po049;
    output po039;
    output po108;
    output po077;
    output po011;
    output po028;
    output po002;
    output po032;
    output po103;
    output po026;
    output po130;
    output po067;
    output po107;
    output po081;
    output po020;
    output po061;
    output po047;
    output po134;
    output po008;
    output po016;
    output po112;
    output po102;
    output po074;
    output po090;
    output po065;
    output po023;
    output po111;
    output po083;
    output po110;
    output po033;
    output po030;
    output po125;
    output po048;
    output po071;
    output po017;
    output po114;
    output po022;
    output po024;
    output po079;
    output po085;
    output po113;
    output po118;
    output po075;
    output po031;
    output po037;
    output po027;
    output po138;
    output po133;
    output po105;
    output po025;
    output po141;
    output po041;
    output po064;
    output po009;
    output po013;
    output po093;
    output po007;
    output po088;
    output po000;
    output po052;
    output po097;
    output po014;
    output po087;
    output po095;
    output po109;
    output po121;
    output po046;
    output po051;
    output po136;
    output po119;
    output po001;
    output po132;
    output po063;
    output po106;
    output po115;
    output po019;

    // Internal wires
    wire not_pi085_8;
    wire not_pi096_4;
    wire and_n788_n1370;
    wire and_n379_not_n1002;
    wire not_n440;
    wire and_pi007_not_n311;
    wire and_not_pi129_2_not_n428;
    wire n945;
    wire and_n704_n1035;
    wire n1247;
    wire and_not_n882_not_n886;
    wire not_pi054_10;
    wire n1570;
    wire and_not_n1470_not_n1471;
    wire n1456;
    wire n1227;
    wire n636;
    wire and_pi073_n958;
    wire not_n1460;
    wire n303;
    wire not_n832;
    wire not_n1271_2;
    wire n351;
    wire and_pi086_not_pi138_403536070;
    wire not_n1472;
    wire not_pi050;
    wire and_pi054_not_n336;
    wire and_not_pi129_10_not_n531;
    wire n1104;
    wire and_not_pi003_3430_n636;
    wire n718;
    wire n1473;
    wire and_not_n1174_not_n1176;
    wire n879;
    wire n410;
    wire n697;
    wire n936;
    wire and_not_pi003_7_n542;
    wire n379;
    wire and_not_n1391_not_n1392;
    wire not_n1552;
    wire and_n385_n697;
    wire and_n754_n755;
    wire n1207;
    wire and_not_pi138_0_n1246;
    wire n613;
    wire and_not_n1285_not_n1287;
    wire and_pi072_not_n1271_1;
    wire and_not_n1187_not_n1189;
    wire n1416;
    wire not_n713;
    wire not_n1492;
    wire and_not_n1218_not_n1220;
    wire not_n1187;
    wire not_n1195;
    wire n1030;
    wire and_n398_n399;
    wire not_pi054;
    wire and_not_pi111_n1621;
    wire and_pi059_not_n1217;
    wire and_n448_n512;
    wire n880;
    wire n1145;
    wire not_n1013;
    wire n873;
    wire n625;
    wire not_pi002_1;
    wire not_pi009_5;
    wire n650;
    wire not_n617;
    wire not_pi026_4;
    wire and_not_pi013_not_pi014;
    wire not_n645;
    wire n1478;
    wire n1540;
    wire and_pi032_not_pi109_1;
    wire n839;
    wire not_n1004;
    wire and_not_pi137_2_not_n1354;
    wire and_n762_not_n777;
    wire not_n575;
    wire not_pi058_7;
    wire and_pi082_not_n409;
    wire and_pi026_pi053;
    wire not_n1215;
    wire n304;
    wire not_n357;
    wire not_n655;
    wire and_not_pi008_n294;
    wire and_pi092_pi106;
    wire not_n1085;
    wire and_not_pi008_3_n449;
    wire n929;
    wire not_pi129_152867006319425761937651857692768264010;
    wire n1245;
    wire and_pi075_not_n1271_4;
    wire not_n1497;
    wire and_pi116_n1578;
    wire not_n1589;
    wire and_not_pi129_725745515342319093317411710931737859674906464051430_not_n1397;
    wire not_pi010_3;
    wire and_pi144_n1386;
    wire and_not_pi041_0_n405;
    wire not_n332;
    wire not_n837;
    wire and_not_n875_not_n879;
    wire and_n705_n1100;
    wire and_pi095_n1324;
    wire not_n1453;
    wire n373;
    wire n362;
    wire not_pi139;
    wire not_n907;
    wire not_n899;
    wire not_n1400;
    wire n656;
    wire n1470;
    wire and_pi057_not_n1194;
    wire and_not_pi129_2824752490_not_n669;
    wire not_n1379;
    wire n1389;
    wire not_pi136_24010;
    wire not_pi044;
    wire not_n1505;
    wire not_n1420;
    wire and_pi093_pi106;
    wire n952;
    wire n1138;
    wire n1414;
    wire and_n777_n790;
    wire not_n870;
    wire and_pi067_not_n1271_0;
    wire and_not_pi015_1_not_n584;
    wire not_n1538;
    wire not_pi007_0;
    wire not_n892;
    wire not_n1150;
    wire n343;
    wire not_n379_9;
    wire not_n624;
    wire not_n1113;
    wire not_pi013_2;
    wire n800;
    wire n748;
    wire and_n420_n421;
    wire not_n1514;
    wire and_pi071_not_n1247_6;
    wire and_not_n654_not_n655;
    wire and_not_n1227_not_n1229;
    wire not_n709;
    wire n384;
    wire po114_driver;
    wire not_n866;
    wire and_not_n965_not_n967;
    wire and_n705_n708;
    wire not_n1271_6;
    wire not_pi056;
    wire po117_driver;
    wire n1095;
    wire and_n445_n480;
    wire not_pi096_1;
    wire not_pi021_0;
    wire n513;
    wire n732;
    wire n811;
    wire and_pi136_not_n1513;
    wire n1340;
    wire and_n401_n698;
    wire not_n379_6;
    wire or_pi129_n1302;
    wire not_n841;
    wire n1459;
    wire n1558;
    wire not_pi053_4;
    wire n1378;
    wire and_pi137_not_n1506;
    wire n571;
    wire and_not_pi024_4_not_pi042_2;
    wire po046_driver;
    wire n604;
    wire not_pi144;
    wire n774;
    wire n593;
    wire not_n919;
    wire and_not_n1000_not_n1003;
    wire not_n979;
    wire not_n1232;
    wire n1413;
    wire not_pi100;
    wire and_pi082_not_n1027;
    wire n831;
    wire not_n1197;
    wire not_n732;
    wire and_n934_n1074;
    wire n1229;
    wire not_n1262;
    wire and_not_pi011_0_not_pi012_1;
    wire not_pi005_0;
    wire and_pi082_not_n645;
    wire po082_driver;
    wire and_n384_n1054;
    wire and_n1251_n1281;
    wire n1609;
    wire n1339;
    wire not_pi003_2824752490;
    wire and_not_pi129_8272697060641711598380789001840137510382698418573894642080092744490_not_n1616;
    wire not_n885;
    wire n971;
    wire po056_driver;
    wire n1342;
    wire not_n696;
    wire and_not_pi096_n714;
    wire and_not_pi145_0_n1271;
    wire and_pi010_not_pi054_5;
    wire not_n353;
    wire not_n719;
    wire not_pi085_9;
    wire not_pi003_273687473400809163430;
    wire n805;
    wire n365;
    wire not_pi002;
    wire and_pi082_not_n391;
    wire n1155;
    wire not_n1144;
    wire and_pi114_not_pi122;
    wire not_pi058;
    wire and_not_n511_not_n519;
    wire n1603;
    wire n659;
    wire n844;
    wire and_n408_n1088;
    wire and_not_n1181_not_n1183;
    wire and_not_n896_not_n900;
    wire not_pi011_0;
    wire and_not_pi129_968890104070_not_n709;
    wire not_n530;
    wire and_not_pi000_not_n306;
    wire n1241;
    wire not_n1377;
    wire and_not_pi129_185621159210175743024531636712070_not_n1096;
    wire and_not_n1613_not_n1615;
    wire and_not_pi129_24118650322570587750381309043265707027354805885055086420058579430_not_n1597;
    wire not_pi085_1;
    wire not_pi003_24010;
    wire not_n764;
    wire and_not_pi085_8_n787;
    wire n649;
    wire n714;
    wire and_n314_n326;
    wire n574;
    wire n504;
    wire n829;
    wire not_n1446;
    wire not_pi027_70;
    wire n675;
    wire not_pi120;
    wire not_n1349;
    wire n630;
    wire not_n358;
    wire not_pi129_1176490;
    wire po100_driver;
    wire n632;
    wire not_n1181;
    wire not_pi007_6;
    wire and_not_n793_not_n797;
    wire po138_driver;
    wire and_not_pi085_0_not_n732;
    wire n777;
    wire not_n844;
    wire n1296;
    wire n1471;
    wire not_n657;
    wire and_not_pi026_70_pi058;
    wire not_pi009;
    wire not_n1019;
    wire and_pi007_n357;
    wire n1403;
    wire n973;
    wire n1217;
    wire or_pi129_n1274;
    wire and_pi053_not_pi085_2;
    wire not_n1386_4;
    wire and_not_n368_not_n370;
    wire po110_driver;
    wire n565;
    wire n1350;
    wire not_n1108;
    wire and_n549_n1614;
    wire not_pi029_1;
    wire and_not_pi026_3430_not_pi053_7;
    wire n551;
    wire not_n1070;
    wire not_pi019_0;
    wire not_n745;
    wire not_n986;
    wire not_n1247_2;
    wire not_pi110;
    wire not_n1545;
    wire and_not_pi003_1_n470;
    wire n391;
    wire and_pi082_not_n1127;
    wire not_n1229;
    wire and_not_pi137_not_pi138;
    wire and_not_n1326_not_n1327;
    wire and_pi096_pi138;
    wire po073_driver;
    wire and_n408_n927;
    wire not_n1005;
    wire n518;
    wire n336;
    wire and_not_pi144_n1249;
    wire not_n1455;
    wire not_n1102;
    wire not_n1336;
    wire and_not_pi116_10_not_n1214;
    wire not_n1096;
    wire not_pi003_7;
    wire not_n625;
    wire n1336;
    wire po024_driver;
    wire not_pi017_1;
    wire not_n903;
    wire n1455;
    wire n1365;
    wire not_n1426;
    wire n1457;
    wire not_pi109_4;
    wire and_not_pi129_3445521474652941107197329863323672432479257983579298060008368490_n1592;
    wire n1441;
    wire n925;
    wire not_n781;
    wire n1200;
    wire n1585;
    wire not_n821;
    wire not_n1121;
    wire not_pi003_8235430;
    wire po062_driver;
    wire not_pi016_2;
    wire not_pi054_9;
    wire not_pi003_138412872010;
    wire and_pi062_n1091;
    wire not_n1169;
    wire and_not_pi043_0_n407;
    wire not_pi027_7;
    wire not_n1076;
    wire not_pi115;
    wire and_not_n379_9_not_n1038;
    wire not_pi129_93874803376477543056490;
    wire n851;
    wire and_not_pi051_1_pi109;
    wire and_n927_n984;
    wire not_n959;
    wire and_n444_n445;
    wire and_not_pi046_1_n388;
    wire and_not_pi009_1_not_pi014_3;
    wire n1075;
    wire po086_driver;
    wire not_n829;
    wire not_n302;
    wire not_pi042_1;
    wire and_not_pi137_8_not_n1519;
    wire not_n328;
    wire n654;
    wire n461;
    wire n854;
    wire and_not_pi002_2_not_pi048_2;
    wire not_n1285;
    wire n1041;
    wire n1071;
    wire and_not_pi141_0_n1271;
    wire and_pi082_not_n692;
    wire n683;
    wire n419;
    wire n1564;
    wire and_not_pi074_not_pi136_9;
    wire not_n1476;
    wire and_not_n1316_not_n1317;
    wire n1502;
    wire and_n354_n373;
    wire and_not_pi043_3_not_n1004;
    wire and_not_pi141_n1249;
    wire n835;
    wire not_pi116_7;
    wire and_n441_n443;
    wire n1191;
    wire and_n583_n587;
    wire n564;
    wire and_pi020_not_n653;
    wire n954;
    wire and_n754_n1154;
    wire and_not_n737_n795;
    wire and_n1583_n1588;
    wire n1171;
    wire and_pi053_not_pi058_4;
    wire and_not_pi142_n1249;
    wire not_n1184;
    wire n890;
    wire n1318;
    wire and_not_pi003_4_n509;
    wire n293;
    wire n321;
    wire n590;
    wire and_pi089_pi138;
    wire not_n1397;
    wire n1017;
    wire n528;
    wire not_n1432;
    wire n966;
    wire not_pi129_8272697060641711598380789001840137510382698418573894642080092744490;
    wire not_pi002_4;
    wire n747;
    wire not_pi053;
    wire not_pi129_797922662976120010;
    wire not_pi146_0;
    wire not_pi070_0;
    wire not_pi138_3430;
    wire and_pi082_not_n920;
    wire and_pi081_pi120;
    wire not_pi026_490;
    wire n1228;
    wire not_pi136_403536070;
    wire not_n1365;
    wire not_pi007_9;
    wire n1064;
    wire not_n1452;
    wire n459;
    wire not_pi123;
    wire n460;
    wire and_n571_n574;
    wire n1581;
    wire not_n930;
    wire n1080;
    wire n941;
    wire not_n1580;
    wire n755;
    wire not_n1225;
    wire and_not_n1503_not_n1507;
    wire n610;
    wire n454;
    wire and_n297_n304;
    wire and_not_pi003_9_n566;
    wire not_n407;
    wire not_n880;
    wire and_pi142_n1414;
    wire and_pi023_pi138;
    wire and_not_pi012_3_n449;
    wire n332;
    wire n352;
    wire n870;
    wire not_n1114;
    wire and_not_n691_not_n694;
    wire not_n869;
    wire and_n407_n580;
    wire po111_driver;
    wire n308;
    wire not_n753;
    wire not_n1366;
    wire and_not_n869_not_n870;
    wire n1208;
    wire and_not_pi044_3_n379;
    wire not_n1414;
    wire not_pi006_2;
    wire not_pi003_8;
    wire n381;
    wire n761;
    wire n905;
    wire and_pi094_not_n1414;
    wire and_not_n959_n962;
    wire not_pi003_0;
    wire n394;
    wire n591;
    wire n1237;
    wire and_not_n379_168070_not_n1158;
    wire n819;
    wire n1517;
    wire not_pi025;
    wire not_n761;
    wire not_n1531;
    wire and_not_pi137_6_not_n1491;
    wire po108_driver;
    wire and_not_pi038_0_not_pi040_0;
    wire n425;
    wire and_pi138_not_n1498;
    wire n817;
    wire n1388;
    wire and_not_n1458_not_n1462;
    wire not_pi085_6;
    wire and_pi100_not_n716;
    wire not_n498;
    wire n1074;
    wire n1335;
    wire n1608;
    wire not_n1459;
    wire or_not_pi122_2_pi129;
    wire and_not_pi070_n577;
    wire not_n1555;
    wire not_n469;
    wire and_n1246_not_n1603;
    wire or_n1499_n1509;
    wire not_pi041;
    wire not_pi011_2;
    wire and_not_n1415_not_n1416;
    wire and_pi079_not_n1325_0;
    wire not_pi041_0;
    wire n1463;
    wire not_n1058;
    wire and_n404_n638;
    wire n1550;
    wire n840;
    wire n980;
    wire not_n1530;
    wire n474;
    wire not_pi028_0;
    wire and_not_n379_6_not_n993;
    wire n1604;
    wire po012_driver;
    wire n1387;
    wire not_pi129_57908879424491981188665523012880962572678888930017262494560649211430;
    wire and_not_pi002_0_not_pi020_0;
    wire not_n589;
    wire and_pi029_not_pi116_5;
    wire and_pi035_n1360;
    wire and_not_n995_n997;
    wire n887;
    wire not_n1271_5;
    wire not_pi129_24010;
    wire not_pi027_4;
    wire and_pi082_not_n956;
    wire not_pi047;
    wire not_pi014;
    wire not_pi129_103677930763188441902487387275962551382129494864490;
    wire n1267;
    wire not_n397;
    wire and_pi137_not_n1487;
    wire n1114;
    wire n960;
    wire n959;
    wire not_n1260;
    wire and_not_n1265_not_n1267;
    wire not_n1475;
    wire not_pi085;
    wire not_pi011_5;
    wire not_n1325_1;
    wire n1338;
    wire n855;
    wire and_n570_n579;
    wire and_not_n1144_not_n1147;
    wire not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490;
    wire and_n399_n568;
    wire n516;
    wire and_not_pi129_3430_not_n565;
    wire and_n380_n688;
    wire and_n379_not_n1122;
    wire n411;
    wire and_not_n911_not_n912;
    wire n1266;
    wire and_not_pi042_not_pi044;
    wire and_not_n1199_not_n1201;
    wire and_pi013_not_pi054_8;
    wire and_n547_n552;
    wire not_n694;
    wire and_n388_n641;
    wire not_pi129_205005145156954906122290109080958673914396262484637238056070;
    wire not_pi069;
    wire n1133;
    wire not_n871;
    wire not_pi129_70316764788835532799945507414768825152637918032230572653232010;
    wire and_pi136_not_pi137_0;
    wire n1268;
    wire n301;
    wire not_pi044_0;
    wire and_not_n1334_not_n1335;
    wire n1059;
    wire and_pi075_n1057;
    wire not_pi138_1;
    wire n1582;
    wire n807;
    wire and_n1251_n1256;
    wire not_n1417;
    wire and_n640_n644;
    wire not_n367;
    wire and_not_pi061_not_pi118;
    wire n1201;
    wire n1530;
    wire n713;
    wire not_n1566;
    wire and_not_pi008_0_not_pi021_0;
    wire not_pi100_0;
    wire n1092;
    wire n772;
    wire n1409;
    wire not_n395;
    wire not_pi136_57648010;
    wire not_pi047_3;
    wire not_n1130;
    wire and_not_pi140_0_n1271;
    wire and_not_pi129_19773267430_not_n682;
    wire n550;
    wire and_not_pi026_490_pi037;
    wire and_not_n1565_not_n1566;
    wire n852;
    wire and_n976_n978;
    wire not_n780;
    wire and_n312_n357;
    wire and_not_n1295_not_n1297;
    wire and_not_pi072_not_pi138_2;
    wire po087_driver;
    wire and_not_pi003_57648010_n785;
    wire and_n927_n991;
    wire n1220;
    wire not_pi129_1181813865805958799768684143120019644340385488367699234582870392070;
    wire not_n1064;
    wire not_pi020;
    wire n467;
    wire and_not_pi018_1_not_pi021_2;
    wire and_n294_n355;
    wire and_not_pi003_16284135979104490_n1532;
    wire and_not_pi106_9_not_n943_0;
    wire not_n662;
    wire not_pi129_225393402906922580878632490;
    wire not_pi129_6;
    wire n769;
    wire not_n968;
    wire n1010;
    wire and_n381_n387;
    wire not_n379_3430;
    wire n1214;
    wire not_pi138_8235430;
    wire n1436;
    wire n530;
    wire n681;
    wire not_n879;
    wire and_not_n1320_not_n1321;
    wire and_not_n1029_not_n1032;
    wire n782;
    wire not_n972;
    wire and_not_n620_not_n624;
    wire n988;
    wire not_n739;
    wire po034_driver;
    wire n1514;
    wire not_n1391;
    wire and_not_pi067_not_pi138_57648010;
    wire and_not_pi047_0_not_pi048_0;
    wire n949;
    wire and_not_n1150_not_n1151;
    wire n1282;
    wire and_pi137_not_n1567;
    wire and_n677_n679;
    wire not_n1124;
    wire and_not_n1178_not_n1179;
    wire and_not_n1485_not_n1486;
    wire n1277;
    wire not_n701;
    wire and_not_pi041_2_not_n968;
    wire n926;
    wire or_n1484_n1494;
    wire not_n1021;
    wire not_pi129_881247870897231951843937366879128181133112010;
    wire n374;
    wire n555;
    wire n317;
    wire not_pi074;
    wire not_pi126;
    wire not_pi054_3;
    wire n424;
    wire n602;
    wire and_not_pi053_0_pi058;
    wire n765;
    wire not_pi022;
    wire n876;
    wire not_pi010_2;
    wire po007_driver;
    wire n815;
    wire not_n728;
    wire and_n322_n516;
    wire not_n531;
    wire not_n716;
    wire not_n878;
    wire not_n927;
    wire and_not_pi010_0_not_pi022_0;
    wire po080_driver;
    wire and_not_pi129_14811132966169777414641055325137507340304213552070_not_n1389;
    wire not_n604;
    wire or_pi129_n1310;
    wire tie1;
    wire not_pi011_3;
    wire and_not_pi139_0_n1271;
    wire n722;
    wire not_n1378;
    wire and_pi016_not_pi054_10;
    wire n1067;
    wire not_n1436;
    wire n1234;
    wire and_not_pi129_85383234134508499009700170379408027452893070589186688070_not_n1430;
    wire not_n1030;
    wire and_n384_n586;
    wire n666;
    wire not_n1556;
    wire n1221;
    wire not_n1450;
    wire and_not_n1034_n1046;
    wire and_not_n1005_n1015;
    wire not_pi116_8;
    wire and_not_pi001_not_n352;
    wire not_n799;
    wire n1150;
    wire not_n983;
    wire n1511;
    wire not_n363;
    wire and_n385_n698;
    wire n670;
    wire not_n1090;
    wire and_pi082_not_n1055;
    wire n502;
    wire and_pi065_not_n1247_2;
    wire n658;
    wire n1395;
    wire not_pi085_490;
    wire not_pi106_2;
    wire n729;
    wire not_po129;
    wire and_not_pi129_26517308458596534717790233816010_not_n1076;
    wire not_n394;
    wire and_pi044_pi082;
    wire n1442;
    wire n1244;
    wire n865;
    wire or_pi129_pi134;
    wire not_n1280;
    wire and_pi092_not_n1386_3;
    wire po005_driver;
    wire not_pi007_5;
    wire not_n482;
    wire and_n450_n610;
    wire and_pi082_not_n985;
    wire po026_driver;
    wire n357;
    wire not_pi007;
    wire not_n410;
    wire and_n927_n929;
    wire and_not_n940_not_n1136;
    wire po083_driver;
    wire n1021;
    wire n736;
    wire not_n576;
    wire n794;
    wire and_pi074_n932;
    wire and_not_n1349_not_n1353;
    wire and_not_pi010_not_n324;
    wire not_n472;
    wire and_not_pi028_0_n548;
    wire not_n1173;
    wire n1298;
    wire n1081;
    wire not_pi110_5;
    wire not_n1405;
    wire n693;
    wire n1072;
    wire n382;
    wire and_not_pi085_6_not_n849;
    wire n994;
    wire n620;
    wire and_pi054_not_pi059_0;
    wire not_n922;
    wire po113_driver;
    wire and_not_n379_5_not_n973;
    wire and_n918_n1043;
    wire not_pi003_6782230728490;
    wire not_n1308;
    wire n969;
    wire and_not_n969_n981;
    wire n294;
    wire and_n1087_n1120;
    wire not_pi058_0;
    wire n1596;
    wire not_pi116_3;
    wire not_n884;
    wire not_n379_10;
    wire and_pi063_not_n1247_0;
    wire n1487;
    wire n315;
    wire not_n794_0;
    wire n430;
    wire not_n1471;
    wire and_n419_n473;
    wire n801;
    wire not_n1596;
    wire not_n311;
    wire not_n656;
    wire not_n908;
    wire and_not_n425_not_n427;
    wire not_pi069_0;
    wire or_pi123_pi129;
    wire and_n536_n537;
    wire and_pi030_not_pi109;
    wire and_pi082_not_n949;
    wire not_pi138_70;
    wire n579;
    wire n1314;
    wire n1358;
    wire n542;
    wire not_n742;
    wire not_pi129_113988951853731430;
    wire and_pi026_pi116;
    wire not_pi095;
    wire and_pi082_not_n394;
    wire n784;
    wire not_n1470;
    wire and_not_pi027_6_not_n804;
    wire and_not_pi136_2824752490_pi140;
    wire not_pi043;
    wire and_not_pi044_0_n401;
    wire not_n861;
    wire po058_driver;
    wire not_pi004_2;
    wire and_not_pi129_168070_not_n601;
    wire not_pi110_6;
    wire and_n383_n384;
    wire not_n795;
    wire and_n404_n406;
    wire n1086;
    wire n1126;
    wire n1182;
    wire and_not_pi129_8_not_n508;
    wire n541;
    wire not_n1344;
    wire and_pi002_n645;
    wire and_n1246_not_n1421;
    wire and_not_pi085_3430_not_n725_0;
    wire po003_driver;
    wire and_pi033_pi109;
    wire n1505;
    wire n323;
    wire n492;
    wire not_pi026_70;
    wire and_pi008_not_pi054_3;
    wire and_not_pi040_2_not_n952;
    wire not_n391;
    wire not_n914;
    wire n1602;
    wire and_not_pi022_3_n449;
    wire n685;
    wire n810;
    wire n449;
    wire not_pi109;
    wire n409;
    wire n1084;
    wire not_n333;
    wire and_not_pi010_2_pi022;
    wire and_n927_n1126;
    wire n1568;
    wire not_n1127;
    wire po019_driver;
    wire not_n845;
    wire n1205;
    wire not_n653;
    wire and_pi035_not_pi109_4;
    wire n742;
    wire n299;
    wire and_n814_n1169;
    wire and_not_pi050_2_n391;
    wire n951;
    wire n469;
    wire not_pi045_2;
    wire po102_driver;
    wire and_not_pi003_1176490_n759;
    wire not_n840;
    wire not_pi109_0;
    wire n499;
    wire and_n638_n1110;
    wire and_not_pi129_1176490_not_n617;
    wire and_n934_n1094;
    wire not_n634;
    wire not_pi043_0;
    wire n1589;
    wire not_pi027_3;
    wire not_n1271_0;
    wire n1044;
    wire not_pi003_2;
    wire or_pi129_n1322;
    wire and_not_n472_not_n482;
    wire and_n490_n492;
    wire and_not_n350_n351;
    wire and_n381_n406;
    wire n405;
    wire n1371;
    wire not_pi041_1;
    wire n417;
    wire and_pi033_pi136;
    wire n746;
    wire n566;
    wire n1222;
    wire n1451;
    wire and_pi145_n1414;
    wire not_pi039_0;
    wire n1238;
    wire not_n1271_4;
    wire not_n792;
    wire not_n1478;
    wire not_n1265;
    wire n1467;
    wire n331;
    wire n768;
    wire n1301;
    wire n1353;
    wire not_n737;
    wire n617;
    wire n1096;
    wire not_pi054_0;
    wire n773;
    wire n776;
    wire not_pi008_2;
    wire po037_driver;
    wire n745;
    wire and_pi006_not_pi012_4;
    wire and_n1246_not_n1585;
    wire and_pi137_not_n1362;
    wire n1065;
    wire and_not_pi143_0_n1249;
    wire and_not_pi014_2_pi054;
    wire not_n915;
    wire n1042;
    wire po103_driver;
    wire n837;
    wire n1121;
    wire not_n1615;
    wire not_n1191;
    wire n892;
    wire n1561;
    wire po094_driver;
    wire and_not_pi129_11044276742439206463052992010_not_n1013;
    wire n1223;
    wire and_not_pi071_n647;
    wire not_n1233;
    wire not_n858;
    wire n396;
    wire n453;
    wire n1033;
    wire and_not_n836_not_n840;
    wire and_not_pi013_1_pi014;
    wire n588;
    wire n1559;
    wire not_n726_0;
    wire not_n853;
    wire not_pi109_1;
    wire and_n379_not_n1065;
    wire n1165;
    wire and_not_pi122_1_n1240;
    wire not_pi113_0;
    wire n1109;
    wire not_pi110_7;
    wire n1190;
    wire n383;
    wire and_n1192_n1196;
    wire or_n1355_n1363;
    wire n1513;
    wire and_pi093_not_n1386_4;
    wire n940;
    wire and_not_pi011_3_n449;
    wire and_not_n1215_not_n1216;
    wire n1575;
    wire n1325;
    wire and_not_n1395_not_n1396;
    wire not_pi129_1577753820348458066150427430;
    wire not_pi017_2;
    wire and_pi145_n1325;
    wire n597;
    wire n720;
    wire not_pi122_2;
    wire not_n508;
    wire not_pi045_3;
    wire n1327;
    wire n1360;
    wire not_pi138_57648010;
    wire not_n1441;
    wire and_n728_n737;
    wire and_not_n1555_not_n1559;
    wire n1554;
    wire n490;
    wire and_pi097_pi138;
    wire n327;
    wire n1381;
    wire and_not_n721_not_n733;
    wire n738;
    wire not_n1525;
    wire n1005;
    wire n822;
    wire n953;
    wire not_pi129_168070;
    wire n1090;
    wire and_not_pi129_12197604876358357001385738625629718207556152941312384010_not_n1426;
    wire and_n344_n374;
    wire and_n448_n491;
    wire not_pi025_1;
    wire n1230;
    wire not_n338;
    wire and_not_pi129_29286449308136415160327158440136953416342323212091034008010_not_n1442;
    wire n1461;
    wire n1488;
    wire and_pi081_not_pi138_1176490;
    wire po059_driver;
    wire not_pi008_1;
    wire po133_driver;
    wire not_pi003_1176490;
    wire and_not_pi047_3_not_n1067;
    wire not_pi018_1;
    wire not_n891;
    wire and_n404_n970;
    wire n942;
    wire n992;
    wire n1320;
    wire and_not_n1601_not_n1602;
    wire and_n355_n488;
    wire not_pi122;
    wire n624;
    wire and_n573_n689;
    wire and_not_n924_n938;
    wire and_not_pi018_not_pi019;
    wire not_n798;
    wire and_not_pi085_9_not_n1188;
    wire n1243;
    wire or_pi129_n1306;
    wire not_n757;
    wire and_not_pi126_pi132;
    wire not_pi022_4;
    wire n456;
    wire and_n344_n416;
    wire and_pi037_not_pi109_6;
    wire n586;
    wire not_pi028;
    wire and_pi086_not_n1325_5;
    wire and_pi054_n1610;
    wire po119_driver;
    wire not_n1404;
    wire po141_driver;
    wire and_pi036_pi109;
    wire and_pi060_pi109;
    wire not_n573;
    wire n1068;
    wire and_not_pi045_not_pi048;
    wire not_n1300;
    wire and_pi048_n1041;
    wire not_pi009_4;
    wire and_not_pi075_not_pi138_490;
    wire n553;
    wire and_not_n1119_not_n1123;
    wire not_pi005;
    wire n1460;
    wire and_not_n779_not_n780;
    wire n1493;
    wire and_not_pi003_n438;
    wire n503;
    wire and_n379_not_n1031;
    wire n432;
    wire n1039;
    wire and_not_pi097_1_n755;
    wire and_n382_n385;
    wire n1166;
    wire not_pi129_725745515342319093317411710931737859674906464051430;
    wire n509;
    wire n809;
    wire n1592;
    wire not_n1342;
    wire not_n1358;
    wire n806;
    wire n733;
    wire not_pi136_3430;
    wire and_n1093_n1095;
    wire and_not_pi007_0_pi013;
    wire n646;
    wire n1037;
    wire n1093;
    wire and_n918_n919;
    wire not_n721;
    wire n1631;
    wire and_not_n735_not_n744;
    wire n389;
    wire not_pi116_10;
    wire n1285;
    wire and_n381_n405;
    wire n1088;
    wire not_n1267;
    wire not_n1052;
    wire n752;
    wire n1422;
    wire and_not_pi136_0_pi137;
    wire and_not_pi021_3_pi054;
    wire and_not_n1514_not_n1518;
    wire and_n448_n504;
    wire not_n812;
    wire n489;
    wire n1273;
    wire not_n1629;
    wire not_n1317;
    wire and_not_n523_not_n530;
    wire not_n805;
    wire n369;
    wire and_pi082_not_n1080;
    wire n1179;
    wire n787;
    wire n823;
    wire not_pi137_3;
    wire and_not_n1544_not_n1548;
    wire and_not_pi085_70_n1212;
    wire and_not_pi058_10_n1206;
    wire and_not_pi024_2_not_n695;
    wire n790;
    wire n575;
    wire not_n1217;
    wire and_n359_n361;
    wire and_not_n1428_not_n1429;
    wire not_pi046_1;
    wire not_n777;
    wire po054_driver;
    wire not_pi051_0;
    wire not_pi021_1;
    wire and_not_pi024_0_not_pi045_0;
    wire n576;
    wire and_n356_n372;
    wire n1386;
    wire not_pi003;
    wire and_not_pi129_490_not_n554;
    wire n614;
    wire n1408;
    wire and_n748_n756;
    wire n465;
    wire n326;
    wire and_not_pi097_n724;
    wire not_n315;
    wire n781;
    wire n878;
    wire and_not_pi129_77309937197074445241370944070_not_n983_0;
    wire n633;
    wire and_n649_n651;
    wire n648;
    wire n1202;
    wire not_n725_0;
    wire not_n1424;
    wire and_not_pi014_1_n347;
    wire and_not_pi025_1_not_pi028_1;
    wire and_pi098_pi106;
    wire n452;
    wire and_not_pi129_1070069044235980333563563003849377848070_not_n1209;
    wire not_n1421_2;
    wire and_n787_n847;
    wire and_pi145_n1386;
    wire and_n448_n545;
    wire not_n1321;
    wire not_pi100_2;
    wire and_not_pi003_490_n626;
    wire n704;
    wire n1370;
    wire not_pi129_248930711762415449007872216849586085868492917169640490;
    wire n402;
    wire not_n1515;
    wire or_n1469_n1479;
    wire and_n369_n431;
    wire or_pi129_n1283;
    wire n912;
    wire po053_driver;
    wire not_pi014_3;
    wire n672;
    wire not_pi027_0;
    wire n1106;
    wire not_n379_24010;
    wire n1152;
    wire n1189;
    wire n1385;
    wire not_n1522;
    wire and_not_pi129_1435036016098684342856030763566710717400773837392460666392490_not_n1531;
    wire and_not_pi129_57908879424491981188665523012880962572678888930017262494560649211430_not_n724;
    wire and_not_pi003_10_n602;
    wire and_not_pi085_5_not_n808;
    wire and_not_pi044_1_pi082;
    wire and_not_n1104_n1116;
    wire n370;
    wire n1586;
    wire n1257;
    wire not_pi137_8;
    wire n1496;
    wire not_pi054_8;
    wire not_pi136_2824752490;
    wire and_n1223_n1224;
    wire not_pi058_6;
    wire not_n1466;
    wire not_pi045_0;
    wire not_n947;
    wire not_n1000;
    wire and_not_n1556_not_n1557;
    wire and_pi074_not_n1271_3;
    wire not_n826;
    wire and_n515_n517;
    wire n324;
    wire n407;
    wire n443;
    wire and_not_n1276_not_n1277;
    wire not_pi066;
    wire not_n1188;
    wire and_n638_n928;
    wire not_n923;
    wire not_pi010_1;
    wire not_n1107;
    wire n1425;
    wire and_n369_n528;
    wire and_n473_n474;
    wire and_not_n1424_not_n1425;
    wire n605;
    wire n1098;
    wire and_not_pi007_6_n449;
    wire and_not_pi002_1_not_pi045_3;
    wire n609;
    wire n1521;
    wire and_not_pi145_n1249;
    wire n418;
    wire n780;
    wire not_pi141_0;
    wire and_pi096_n1370;
    wire n1103;
    wire not_n703;
    wire and_not_pi136_8235430_not_n1564;
    wire not_n758;
    wire n694;
    wire n1444;
    wire not_pi146;
    wire and_not_n696_n711;
    wire n1031;
    wire n598;
    wire po129_driver;
    wire po006_driver;
    wire n519;
    wire n1260;
    wire and_n402_n408;
    wire not_pi039;
    wire and_not_n1081_not_n1083;
    wire not_n1559;
    wire and_not_pi106_1_not_n878;
    wire n726;
    wire not_n1423;
    wire not_pi049_0;
    wire n1169;
    wire n628;
    wire n447;
    wire not_pi085_0;
    wire not_n1040;
    wire n1454;
    wire n1468;
    wire and_not_pi068_pi136;
    wire not_n1564;
    wire n339;
    wire n967;
    wire and_pi082_not_n573;
    wire not_n1485;
    wire not_n1247_6;
    wire and_not_pi096_2_n830;
    wire and_n448_n535;
    wire not_pi002_2;
    wire and_n538_n539;
    wire and_not_n578_n592;
    wire not_pi007_2;
    wire and_n1054_n1059;
    wire po109_driver;
    wire and_pi125_pi138;
    wire and_pi116_n737;
    wire not_n336;
    wire and_not_n837_not_n838;
    wire not_n941;
    wire not_pi009_6;
    wire n1304;
    wire not_pi010_0;
    wire not_n943_0;
    wire n1215;
    wire and_not_n486_not_n494;
    wire not_pi100_1;
    wire and_pi032_pi109;
    wire not_n591;
    wire not_n1423_0;
    wire and_n380_n1111;
    wire and_n1581_n1583;
    wire not_pi129_125892552985318850263419623839875454447587430;
    wire n669;
    wire not_n320;
    wire n663;
    wire po051_driver;
    wire n1046;
    wire po127_driver;
    wire not_pi006_1;
    wire not_pi110_0;
    wire n1020;
    wire and_not_pi003_797922662976120010_n1577;
    wire not_pi040_2;
    wire not_n993;
    wire not_n1123;
    wire not_n685;
    wire and_pi005_not_n332;
    wire not_pi047_4;
    wire and_not_n379_not_n395;
    wire n1506;
    wire not_pi022_2;
    wire not_pi129_6168735096280623662907561568153897267931784070;
    wire n642;
    wire and_n380_n381;
    wire not_pi129_367033682172941254412302110320336601888010;
    wire not_n752;
    wire n1501;
    wire not_n796;
    wire not_pi026_168070;
    wire n494;
    wire n1464;
    wire not_n808;
    wire and_pi085_n718;
    wire and_not_n854_not_n857;
    wire not_pi138_8;
    wire not_n1023;
    wire not_n985;
    wire and_not_n868_not_n872;
    wire not_n1430;
    wire not_n723;
    wire n1236;
    wire not_n1290;
    wire and_not_pi136_3_n1411;
    wire po001_driver;
    wire and_not_pi007_2_not_pi013_2;
    wire not_pi003_3;
    wire and_pi082_not_n992;
    wire n1328;
    wire and_pi096_n1219;
    wire and_pi143_n1386;
    wire n1573;
    wire not_pi042_0;
    wire not_n1354;
    wire n757;
    wire and_not_pi085_7_not_n1177;
    wire n585;
    wire and_not_n1260_not_n1262;
    wire n889;
    wire and_not_n1488_not_n1492;
    wire not_pi003_39098210485829880490;
    wire not_n1542;
    wire po027_driver;
    wire and_not_n1140_n1141;
    wire or_pi129_pi135;
    wire not_pi110_2;
    wire not_n740;
    wire n922;
    wire not_n1216;
    wire and_not_pi129_797922662976120010_not_n873;
    wire n495;
    wire and_not_pi129_2326305139872070_not_n826;
    wire n1177;
    wire and_pi142_n1325;
    wire and_not_pi006_2_n450;
    wire not_pi009_0;
    wire and_n345_n346;
    wire and_n813_n814;
    wire and_pi077_n1009;
    wire n1024;
    wire n814;
    wire n1062;
    wire not_pi085_70;
    wire not_pi067;
    wire n320;
    wire n334;
    wire and_pi038_n641;
    wire n989;
    wire n380;
    wire n607;
    wire and_n560_n563;
    wire not_n660;
    wire n996;
    wire and_pi138_not_n1483;
    wire n481;
    wire n1614;
    wire not_pi027_10;
    wire and_not_pi041_not_pi046;
    wire not_n1248;
    wire n846;
    wire po040_driver;
    wire and_not_n1381_not_n1382;
    wire and_pi093_pi138;
    wire n441;
    wire and_n688_n927;
    wire not_n1425;
    wire and_not_pi009_3_not_pi022_2;
    wire and_not_pi003_3_n496;
    wire n696;
    wire and_not_n713_not_n715;
    wire n298;
    wire and_n723_n727;
    wire not_pi144_0;
    wire and_not_pi004_0_not_pi019_0;
    wire not_n1359;
    wire not_pi058_4;
    wire po090_driver;
    wire n526;
    wire n292;
    wire n545;
    wire or_pi003_not_n377;
    wire and_not_pi042_1_not_n988;
    wire and_not_pi138_8_not_n1478;
    wire n987;
    wire and_not_pi137_7_not_n1502;
    wire n375;
    wire n367;
    wire n1176;
    wire n1052;
    wire not_n301;
    wire not_n454;
    wire n679;
    wire and_not_n1280_not_n1282;
    wire and_not_pi110_0_not_n725;
    wire and_not_pi106_3_not_n892;
    wire n877;
    wire not_n843;
    wire and_pi066_not_n1271;
    wire n1181;
    wire n483;
    wire not_n723_0;
    wire and_pi027_n768;
    wire n923;
    wire not_pi097_0;
    wire n1619;
    wire n1518;
    wire n1193;
    wire n638;
    wire not_n1350;
    wire not_pi138_24010;
    wire n1343;
    wire not_pi007_10;
    wire and_not_pi027_4_n737;
    wire and_not_pi129_597682638941559493067901192655856192170251494124306816490_not_n1434;
    wire not_n428;
    wire not_pi027_9;
    wire not_n862;
    wire not_pi045_4;
    wire and_not_pi129_1577753820348458066150427430_not_n996;
    wire n1432;
    wire n413;
    wire n950;
    wire n997;
    wire po039_driver;
    wire and_not_pi015_not_pi020;
    wire not_pi106_1;
    wire not_n1001;
    wire n1565;
    wire n883;
    wire not_n1044;
    wire n1354;
    wire and_not_pi066_not_pi136_7;
    wire n908;
    wire and_n1251_n1266;
    wire not_n1158;
    wire and_pi140_n1386;
    wire and_pi066_n1129;
    wire po093_driver;
    wire not_n833;
    wire and_pi144_n1325;
    wire and_not_pi003_5_n521;
    wire and_n300_n342;
    wire not_n857;
    wire not_n1032;
    wire and_pi082_not_n404;
    wire not_pi136_1;
    wire not_pi137_9;
    wire not_n1548;
    wire n354;
    wire and_not_pi076_not_pi138_168070;
    wire n1188;
    wire not_pi053_5;
    wire and_n605_n607;
    wire and_not_pi004_not_pi016;
    wire n1504;
    wire n559;
    wire n753;
    wire not_n1292;
    wire n1048;
    wire not_n1084;
    wire n1212;
    wire and_not_pi110_6_n1419;
    wire and_not_pi043_not_pi047;
    wire not_n1297;
    wire n1258;
    wire not_pi045_1;
    wire not_n992;
    wire and_n640_n652;
    wire n711;
    wire and_not_pi050_3_n404;
    wire not_n1603;
    wire not_n319;
    wire and_not_pi110_2_n800;
    wire n863;
    wire n660;
    wire not_pi014_2;
    wire n309;
    wire and_not_pi053_2_not_pi058_1;
    wire and_pi085_n787;
    wire and_not_pi136_1_not_n1352;
    wire not_n690;
    wire not_pi096_0;
    wire and_n502_n506;
    wire n560;
    wire and_not_n1330_not_n1331;
    wire and_not_n1338_not_n1339;
    wire not_pi048_1;
    wire and_not_pi006_0_not_pi012_0;
    wire n621;
    wire not_pi143_0;
    wire not_pi136_8;
    wire not_pi106_6;
    wire n1027;
    wire and_not_n1448_not_n1449;
    wire and_n487_n623;
    wire and_pi026_n718;
    wire or_pi129_n1314;
    wire n442;
    wire n444;
    wire not_n755;
    wire not_pi117;
    wire n1141;
    wire and_not_n1290_not_n1292;
    wire not_pi002_0;
    wire n1073;
    wire not_pi003_2326305139872070;
    wire not_n733;
    wire not_n1549;
    wire not_pi008;
    wire and_not_n353_not_n375;
    wire n961;
    wire and_not_n829_not_n834;
    wire and_not_n1255_not_n1257;
    wire and_pi138_n1412;
    wire not_pi129_10045252112690790399992215344966975021805416861747224664747430;
    wire not_pi011_6;
    wire n1132;
    wire and_not_pi106_4_not_n899;
    wire not_n873;
    wire n464;
    wire n1094;
    wire not_pi026_9;
    wire n1043;
    wire not_n1541;
    wire not_pi129_302268019717750559482470516839540966128657419430;
    wire not_pi136_7;
    wire and_pi082_not_n927;
    wire and_pi082_not_n919;
    wire n1591;
    wire and_n379_not_n1050;
    wire not_n1602;
    wire and_n1606_n1607;
    wire po115_driver;
    wire n657;
    wire and_pi045_n1041;
    wire n1003;
    wire n1053;
    wire po126_driver;
    wire not_n1388;
    wire n1283;
    wire n1149;
    wire not_pi052;
    wire not_pi048_2;
    wire and_pi095_not_n1423;
    wire and_pi137_not_n1463;
    wire not_n413;
    wire and_not_pi048_3_not_n1084;
    wire not_n327;
    wire and_not_pi028_n460;
    wire n537;
    wire n783;
    wire and_not_pi026_6_not_pi100_1;
    wire n857;
    wire n640;
    wire and_not_n379_2_not_n701;
    wire not_n770;
    wire and_not_pi100_2_pi116;
    wire and_pi082_not_n930;
    wire n1580;
    wire n1453;
    wire not_n950;
    wire not_n905;
    wire not_n1072;
    wire and_not_n876_not_n877;
    wire not_n1214;
    wire not_n1361;
    wire n1022;
    wire n527;
    wire and_pi019_not_pi054_3430;
    wire not_pi096;
    wire not_n379_4;
    wire not_n1053;
    wire and_pi037_n1360;
    wire not_n1540;
    wire not_n796_0;
    wire n1218;
    wire not_n898;
    wire n918;
    wire n701;
    wire and_not_pi017_1_pi054;
    wire not_pi044_2;
    wire not_n1048;
    wire n1116;
    wire and_n503_n525;
    wire not_n339;
    wire and_not_pi053_8_n1211;
    wire and_pi087_not_pi138_3;
    wire and_not_pi003_19773267430_n1153;
    wire not_n314;
    wire n1407;
    wire not_pi050_3;
    wire not_pi129_8;
    wire and_n1251_n1324;
    wire po042_driver;
    wire and_not_pi116_0_n747;
    wire n1158;
    wire or_pi129_n1258;
    wire not_n975;
    wire not_n379_70;
    wire n1379;
    wire not_pi096_2;
    wire and_not_n740_not_n741;
    wire not_n1183;
    wire and_not_n1511_not_n1512;
    wire and_pi026_not_pi027_5;
    wire and_n638_n954;
    wire not_n379;
    wire not_n1474;
    wire not_n1174;
    wire and_not_pi129_13410686196639649008070_not_n908;
    wire not_n987;
    wire n653;
    wire n1137;
    wire and_pi057_not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490;
    wire not_n806;
    wire not_pi000;
    wire and_n357_n549;
    wire and_pi026_not_pi058_6;
    wire not_n635;
    wire n1524;
    wire and_not_n790_not_n791;
    wire n665;
    wire and_not_pi058_7_n1175;
    wire n1549;
    wire and_n776_n801;
    wire and_not_pi129_2115876138024253916377293617876786762900601936010_not_n1383;
    wire not_pi054_1176490;
    wire not_pi016_1;
    wire and_not_pi044_2_n649;
    wire not_n1282;
    wire and_n344_n348;
    wire po014_driver;
    wire n505;
    wire n1008;
    wire and_pi049_n411;
    wire and_n314_n322;
    wire n387;
    wire not_pi005_5;
    wire not_n834;
    wire po095_driver;
    wire n1198;
    wire n1001;
    wire not_n668;
    wire n482;
    wire n1097;
    wire n1344;
    wire not_pi129_47475615099430;
    wire and_not_pi004_1_not_pi018_3;
    wire not_n1486;
    wire po013_driver;
    wire n1560;
    wire not_pi024_1;
    wire n920;
    wire and_not_pi129_5585458640832840070_not_n880;
    wire not_pi129_32199057558131797268376070;
    wire and_n332_n500;
    wire not_n1226;
    wire not_pi007_3;
    wire n1584;
    wire n1272;
    wire po000_driver;
    wire n1112;
    wire and_pi146_n1386;
    wire not_n1449;
    wire not_n765;
    wire and_pi082_not_n1325_3;
    wire n1069;
    wire and_pi082_not_n575;
    wire not_n1616;
    wire and_pi082_not_n1113;
    wire n734;
    wire n799;
    wire not_pi049_1;
    wire and_pi082_not_n1121;
    wire n739;
    wire n727;
    wire n834;
    wire and_not_pi005_5_n596;
    wire and_n401_n926;
    wire not_n1506;
    wire n345;
    wire and_not_n1312_not_n1313;
    wire and_not_pi026_0_not_pi085_1;
    wire not_pi129_273687473400809163430;
    wire not_pi072;
    wire n1566;
    wire n866;
    wire and_not_pi085_not_pi110;
    wire and_not_n864_not_n865;
    wire or_pi129_n1318;
    wire n962;
    wire and_n390_n977;
    wire n360;
    wire or_pi129_n1288;
    wire n476;
    wire and_not_n362_not_n363;
    wire and_n293_n296;
    wire n932;
    wire and_not_n1300_not_n1301;
    wire not_n370;
    wire not_n1038;
    wire and_not_n726_1_n787;
    wire n1274;
    wire n1206;
    wire n325;
    wire n393;
    wire and_not_pi058_8_not_n1190;
    wire n1028;
    wire and_not_pi026_168070_n1375;
    wire not_n1473;
    wire not_pi013_1;
    wire n297;
    wire not_pi109_3;
    wire n1127;
    wire not_pi026_24010;
    wire and_not_n582_not_n588;
    wire po076_driver;
    wire and_not_pi129_52433383167563036344614587188619514555430_n1241;
    wire n1397;
    wire not_n1092;
    wire n691;
    wire and_not_pi129_0_not_n376;
    wire and_not_pi129_8235430_not_n625;
    wire n1004;
    wire not_pi129_2;
    wire not_pi054_6;
    wire not_n584;
    wire and_pi046_pi082;
    wire n1306;
    wire and_n408_n699;
    wire not_pi136_9;
    wire n991;
    wire not_n731;
    wire not_n882;
    wire and_pi042_n934;
    wire and_not_n1020_not_n1021;
    wire not_pi129_24118650322570587750381309043265707027354805885055086420058579430;
    wire po122_driver;
    wire po030_driver;
    wire not_pi018_0;
    wire not_pi129_138412872010;
    wire and_not_pi110_7_not_pi120;
    wire n1136;
    wire not_n1565;
    wire not_pi047_0;
    wire not_pi014_0;
    wire not_pi129_445676403263631959001900459745680070;
    wire and_not_n1459_not_n1460;
    wire not_pi002_3;
    wire n1002;
    wire not_pi003_5585458640832840070;
    wire not_pi054_2;
    wire and_pi010_n291;
    wire n397;
    wire not_n1295;
    wire and_not_n1068_n1078;
    wire n719;
    wire and_not_n1489_not_n1490;
    wire n1383;
    wire and_not_n767_not_n769;
    wire n699;
    wire and_pi111_pi138;
    wire not_pi053_6;
    wire n512;
    wire not_n1117;
    wire not_n404;
    wire and_not_pi085_4_not_n738_0;
    wire not_n379_8;
    wire and_not_pi005_1_n332;
    wire n404;
    wire not_n1132;
    wire not_n1437;
    wire not_pi003_332329305696010;
    wire not_n1536;
    wire and_n316_n318;
    wire not_pi012_2;
    wire n1089;
    wire not_pi003_1;
    wire not_pi085_4;
    wire not_n1003;
    wire not_pi043_2;
    wire not_pi007_1;
    wire not_n823;
    wire n893;
    wire and_not_n1023_n1024;
    wire and_pi097_not_pi110_3;
    wire not_pi122_1;
    wire and_n1583_n1600;
    wire po052_driver;
    wire not_n1351;
    wire and_pi088_not_n1386;
    wire and_n786_n788;
    wire n536;
    wire n986;
    wire not_pi026_0;
    wire not_n746;
    wire not_pi013_5;
    wire not_n376;
    wire not_n1055;
    wire and_not_pi082_n379;
    wire not_n1190;
    wire n1357;
    wire po002_driver;
    wire and_pi099_not_n1386_6;
    wire n618;
    wire not_n1456;
    wire n1577;
    wire and_n408_n585;
    wire not_pi115_0;
    wire or_n1561_n1568;
    wire not_n996;
    wire not_n1386_1;
    wire and_not_n1108_not_n1112;
    wire and_pi030_pi109;
    wire and_not_pi007_4_n332;
    wire n1185;
    wire not_n364;
    wire and_n675_n680;
    wire n1110;
    wire and_not_n1169_not_n1171;
    wire n981;
    wire not_n1325_4;
    wire not_pi012_6;
    wire and_not_n662_not_n668;
    wire not_n1570;
    wire and_not_n823_not_n825;
    wire and_not_n1350_not_n1351;
    wire n435;
    wire n1211;
    wire and_n927_n1017;
    wire n1483;
    wire not_pi129_52433383167563036344614587188619514555430;
    wire or_n1543_n1550;
    wire not_pi113;
    wire n507;
    wire n1430;
    wire not_n628;
    wire not_n1051;
    wire not_n1401;
    wire not_n1421_0;
    wire and_pi034_not_pi109_3;
    wire not_n1493;
    wire not_pi026_5;
    wire n601;
    wire n707;
    wire n1312;
    wire and_pi076_n974;
    wire and_pi136_not_n1454;
    wire n376;
    wire n1131;
    wire n1543;
    wire not_pi047_1;
    wire not_n1178;
    wire and_not_n1432_not_n1433;
    wire not_pi048_0;
    wire not_pi051_1;
    wire and_n390_n650;
    wire po120_driver;
    wire and_not_pi040_1_not_pi042_0;
    wire and_not_n703_n710;
    wire and_n1251_n1385;
    wire not_n940_0;
    wire n1396;
    wire n508;
    wire and_pi087_not_n1325_6;
    wire not_n1221;
    wire not_n1194;
    wire and_pi091_n1249;
    wire not_pi082;
    wire n514;
    wire and_not_pi059_n356;
    wire and_pi078_not_pi136_8;
    wire n901;
    wire and_pi131_n1245;
    wire and_n927_n971;
    wire not_pi063;
    wire n1607;
    wire not_pi116_70;
    wire n1538;
    wire and_pi089_pi106;
    wire and_not_n953_n963;
    wire and_not_pi106_8_n1137;
    wire and_not_n810_not_n811;
    wire n1424;
    wire not_n1257;
    wire and_not_n1452_not_n1453;
    wire n1494;
    wire and_not_pi016_0_pi054;
    wire n1278;
    wire po136_driver;
    wire not_n1122;
    wire n1562;
    wire n1066;
    wire and_pi146_n1325;
    wire n612;
    wire n1184;
    wire not_n1157;
    wire not_pi003_797922662976120010;
    wire po044_driver;
    wire and_not_n742_n743;
    wire not_pi129_5585458640832840070;
    wire n668;
    wire n347;
    wire not_pi040_0;
    wire and_pi082_not_n407;
    wire not_n1148;
    wire not_n1591;
    wire not_pi059_0;
    wire not_pi138_0;
    wire n333;
    wire n678;
    wire not_pi058_5;
    wire not_n337;
    wire not_pi052_0;
    wire not_n1271_3;
    wire not_n1560;
    wire n1322;
    wire not_n1483;
    wire and_not_pi027_0_n749;
    wire n1246;
    wire not_n1356;
    wire and_not_pi008_1_not_pi011_1;
    wire not_pi106_5;
    wire po137_driver;
    wire and_pi082_not_pi138_7;
    wire n956;
    wire not_n317;
    wire not_n728_0;
    wire n1174;
    wire and_not_pi003_1915812313805664144010_not_n1628;
    wire and_not_n1048_not_n1051;
    wire not_pi129_1;
    wire not_n1462;
    wire and_pi116_n1573;
    wire not_n802;
    wire not_n1172;
    wire and_not_n1248_not_n1252;
    wire not_n1231;
    wire and_pi136_n1243;
    wire not_n1408;
    wire and_not_pi003_39098210485829880490_n1609;
    wire n948;
    wire and_not_pi003_70_n618;
    wire po064_driver;
    wire and_pi090_pi106;
    wire n1115;
    wire and_pi082_not_n656;
    wire and_not_n1481_not_n1482;
    wire and_not_pi025_not_pi029;
    wire n919;
    wire not_pi129_13410686196639649008070;
    wire n771;
    wire and_not_n1496_not_n1497;
    wire n710;
    wire n406;
    wire and_not_pi054_1176490_not_pi113_0;
    wire and_not_pi002_4_not_pi047_4;
    wire and_not_pi117_not_pi122_0;
    wire not_n1246;
    wire and_not_pi004_2_not_pi012_6;
    wire n540;
    wire n319;
    wire n1392;
    wire not_pi026_10;
    wire not_n377;
    wire n728;
    wire po081_driver;
    wire n466;
    wire and_n291_n292;
    wire n310;
    wire n652;
    wire and_pi008_pi021;
    wire and_n311_n341;
    wire n825;
    wire n934;
    wire and_n1026_n1027;
    wire not_pi003_19773267430;
    wire not_n1273;
    wire not_n890;
    wire and_pi138_n1246;
    wire n1445;
    wire and_not_pi026_not_n720;
    wire and_not_pi136_1176490_not_n1558;
    wire n968;
    wire and_pi006_pi012;
    wire and_pi064_not_n1247_1;
    wire not_n717;
    wire not_n1104;
    wire and_not_pi115_0_not_n1421_2;
    wire not_n1386;
    wire and_not_pi058_2_not_n822;
    wire and_not_n648_n659;
    wire not_n1227;
    wire po033_driver;
    wire n1119;
    wire n957;
    wire not_n1334;
    wire and_not_n1356_not_n1357;
    wire and_not_pi053_4_not_n841;
    wire not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070;
    wire and_not_pi065_n396;
    wire and_pi047_n641;
    wire n903;
    wire not_pi003_5;
    wire n1491;
    wire not_n900;
    wire n371;
    wire not_n1482;
    wire not_pi138_490;
    wire n390;
    wire not_n1395;
    wire not_n1467;
    wire and_not_pi129_39098210485829880490_not_n887;
    wire and_n584_n650;
    wire n983;
    wire n1484;
    wire and_not_pi129_9_not_n520;
    wire not_n973;
    wire not_n875;
    wire n938;
    wire not_pi004_1;
    wire and_not_n1064_not_n1066;
    wire and_not_n809_not_n815;
    wire n1508;
    wire n849;
    wire and_n1049_n1054;
    wire n907;
    wire and_not_pi136_403536070_pi141;
    wire not_n581;
    wire and_n403_n405;
    wire n1290;
    wire and_n856_n1223;
    wire n1355;
    wire n1553;
    wire and_not_pi051_not_pi052;
    wire not_pi097_1;
    wire n1438;
    wire not_pi110_3;
    wire and_pi143_n1325;
    wire not_pi026_8;
    wire not_n1562;
    wire not_pi004_0;
    wire and_n1251_n1296;
    wire not_pi008_3;
    wire and_n1251_n1286;
    wire and_pi097_not_n1423_1;
    wire not_pi027_3430;
    wire n1393;
    wire not_n1371;
    wire n626;
    wire and_not_pi005_4_n479;
    wire and_not_n843_0_not_n1575;
    wire n1000;
    wire not_n1002;
    wire and_pi004_not_pi054;
    wire not_pi007_8;
    wire and_not_n557_not_n564;
    wire n1423;
    wire not_pi129_70;
    wire not_pi015_1;
    wire and_pi008_not_pi017_3;
    wire not_pi018_3;
    wire not_pi027_1;
    wire and_n1086_n1087;
    wire n798;
    wire n328;
    wire n1070;
    wire and_not_pi129_32199057558131797268376070_not_n961;
    wire not_n1320;
    wire not_pi056_0;
    wire not_n437;
    wire and_pi021_not_pi054_24010;
    wire and_pi146_n1414;
    wire n778;
    wire not_n848;
    wire and_n776_n778;
    wire n475;
    wire n549;
    wire n763;
    wire and_n688_n976;
    wire n606;
    wire and_not_pi011_5_n311;
    wire n698;
    wire n1572;
    wire and_pi029_not_pi097_0;
    wire and_not_pi129_1915812313805664144010_not_n901;
    wire not_pi116_4;
    wire n767;
    wire not_n1202;
    wire n361;
    wire and_n369_n417;
    wire and_n417_n598;
    wire n1076;
    wire n1036;
    wire not_n1383;
    wire not_pi027_2;
    wire and_not_pi116_2_not_n796;
    wire and_n927_n955;
    wire n937;
    wire n344;
    wire not_pi129_3;
    wire and_n568_n572;
    wire not_pi015;
    wire and_not_n883_not_n884;
    wire not_pi136_8235430;
    wire and_not_n1085_n1098;
    wire not_n943;
    wire n1197;
    wire n623;
    wire n539;
    wire n1331;
    wire po104_driver;
    wire not_pi005_4;
    wire not_pi136;
    wire n318;
    wire not_pi136_168070;
    wire not_n983_0;
    wire n544;
    wire and_pi141_n1325;
    wire not_n306;
    wire n583;
    wire po112_driver;
    wire not_pi013_0;
    wire n759;
    wire n935;
    wire and_pi100_not_n766;
    wire n1262;
    wire and_n838_n851;
    wire n927;
    wire not_pi129_57648010;
    wire not_n1029;
    wire n1482;
    wire n573;
    wire and_not_pi045_2_n399;
    wire and_not_pi027_not_n734;
    wire po041_driver;
    wire and_not_pi085_490_not_n1221;
    wire n521;
    wire not_pi021;
    wire not_pi085_3430;
    wire and_n819_n820;
    wire n1035;
    wire not_n1140;
    wire n891;
    wire n450;
    wire and_not_pi026_9_not_n853;
    wire not_n948;
    wire and_not_n1580_not_n1584;
    wire and_n663_n666;
    wire not_pi129_4;
    wire not_n600;
    wire and_not_pi129_152867006319425761937651857692768264010_not_n1202;
    wire n645;
    wire and_not_pi085_10_n1187;
    wire and_not_n1534_not_n1535;
    wire and_not_pi003_0_n456;
    wire n1253;
    wire and_not_n799_n807;
    wire and_not_n1195_not_n1197;
    wire and_pi136_not_pi138_4;
    wire and_pi082_not_n690;
    wire not_pi112;
    wire and_not_pi137_9_not_n1542;
    wire not_n1513;
    wire and_pi085_n774;
    wire n1369;
    wire n862;
    wire and_n379_not_n966;
    wire n531;
    wire po128_driver;
    wire n1167;
    wire not_n843_0;
    wire and_pi082_not_n1089;
    wire not_pi038;
    wire and_pi124_pi138;
    wire not_pi038_1;
    wire n312;
    wire and_pi140_n1325;
    wire not_n593;
    wire not_n455;
    wire not_pi054_3430;
    wire and_not_pi129_6168735096280623662907561568153897267931784070_not_n1367;
    wire not_n390;
    wire n1134;
    wire and_not_pi129_445676403263631959001900459745680070_not_n1142;
    wire and_not_pi062_not_pi138_1;
    wire not_pi018;
    wire not_n595;
    wire and_not_pi027_10_not_n1180;
    wire and_n629_n632;
    wire n479;
    wire not_pi029_0;
    wire and_pi070_not_n1247_5;
    wire n1349;
    wire not_pi129_35561530251773635572553173835655155124070416738520070;
    wire n1597;
    wire not_n565;
    wire n1536;
    wire and_n569_n570;
    wire n517;
    wire not_pi085_2;
    wire n1057;
    wire and_not_n846_not_n848;
    wire not_pi012_4;
    wire n1250;
    wire and_not_pi129_225393402906922580878632490_not_n979;
    wire and_pi078_not_n1325;
    wire not_pi116;
    wire n1023;
    wire and_pi032_pi136;
    wire and_not_pi003_6782230728490_n1210;
    wire n314;
    wire and_not_n1164_0_not_n1170;
    wire and_pi002_not_n412;
    wire n915;
    wire not_n782;
    wire not_pi043_3;
    wire and_n487_n667;
    wire n322;
    wire not_pi136_0;
    wire not_n1138;
    wire n1276;
    wire not_pi129_968890104070;
    wire and_not_pi003_113988951853731430_n1572;
    wire not_pi049;
    wire not_pi138_9;
    wire n764;
    wire and_not_n321_not_n323;
    wire and_not_pi115_pi138;
    wire and_not_n1359_not_n1361;
    wire not_pi013_4;
    wire not_n379_0;
    wire not_pi005_2;
    wire not_n313;
    wire and_not_pi129_7_not_n495;
    wire and_pi067_not_n379_8;
    wire n440;
    wire n445;
    wire and_pi097_pi116;
    wire n743;
    wire not_n669;
    wire not_pi129_7;
    wire and_not_pi146_0_n1271;
    wire and_not_pi137_70_pi138;
    wire not_n886;
    wire and_not_pi106_6_not_n913;
    wire and_not_n1436_not_n1437;
    wire n395;
    wire not_n362;
    wire n1026;
    wire not_pi140;
    wire not_n1027;
    wire n1018;
    wire n1085;
    wire and_not_n1072_n1077;
    wire n1168;
    wire not_n738_0;
    wire and_pi058_not_pi116_7;
    wire not_n1176;
    wire and_not_pi003_8235430_n771;
    wire and_pi031_n1360;
    wire and_pi084_not_n1325_4;
    wire not_n1403;
    wire po079_driver;
    wire n1172;
    wire not_n427;
    wire not_pi110_4;
    wire and_n291_n676;
    wire and_pi029_pi110;
    wire not_pi019_1;
    wire not_pi003_47475615099430;
    wire and_pi025_not_n726;
    wire n1224;
    wire not_n1332;
    wire po070_driver;
    wire n741;
    wire n797;
    wire n1019;
    wire po061_driver;
    wire not_n1501;
    wire n635;
    wire not_n601;
    wire not_n436;
    wire not_pi012_3;
    wire not_n933;
    wire and_n389_n948;
    wire not_pi129_77309937197074445241370944070;
    wire and_pi082_not_n408;
    wire and_not_pi129_367033682172941254412302110320336601888010_not_n1328;
    wire not_pi129_10;
    wire n756;
    wire not_pi129_3430;
    wire and_pi031_not_pi109_0;
    wire not_n876;
    wire not_n1018;
    wire n1120;
    wire not_n1595;
    wire not_n411;
    wire not_n1247_4;
    wire not_pi137_10;
    wire not_pi145_0;
    wire not_pi136_490;
    wire n1433;
    wire and_pi082_not_n1001;
    wire n1537;
    wire and_n399_n697;
    wire n577;
    wire n758;
    wire not_n1328;
    wire and_n819_n824;
    wire and_n311_n312;
    wire not_n1037;
    wire not_pi071;
    wire not_pi129_2824752490;
    wire n1056;
    wire not_pi054_70;
    wire not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430;
    wire and_not_n1010_n1014;
    wire po018_driver;
    wire or_pi129_n1253;
    wire n1271;
    wire and_not_n365_not_n366;
    wire n1571;
    wire n1194;
    wire not_n1081;
    wire not_n1338;
    wire n538;
    wire and_n736_n940;
    wire n998;
    wire not_n1511;
    wire not_n917;
    wire n570;
    wire or_pi129_n1278;
    wire not_pi129_9;
    wire not_n423;
    wire not_pi050_2;
    wire not_n1386_6;
    wire and_n448_n476;
    wire not_n1487;
    wire and_not_pi003_2824752490_n859;
    wire and_n391_n572;
    wire and_pi061_n686;
    wire n1180;
    wire not_pi003_16284135979104490;
    wire n1248;
    wire n1615;
    wire and_not_pi129_4183778472590916451475308348590993345191760458870147715430_not_n1438;
    wire not_n715;
    wire and_not_n983_not_n987;
    wire n1544;
    wire and_not_pi136_3430_not_n1523;
    wire and_not_n730_not_n731;
    wire n493;
    wire not_pi003_968890104070;
    wire not_pi003_168070;
    wire and_n642_n643;
    wire n1356;
    wire not_n494;
    wire n1334;
    wire and_not_pi013_3_not_n364;
    wire not_n495;
    wire and_not_pi136_490_not_n1517;
    wire po021_driver;
    wire and_not_n1538_not_n1539;
    wire not_n852;
    wire not_n1389;
    wire not_pi045;
    wire and_not_n534_not_n540;
    wire and_pi136_not_n1348;
    wire not_n1498;
    wire n1078;
    wire not_n335;
    wire n1292;
    wire not_pi026_7;
    wire and_not_pi112_n1324;
    wire not_n648;
    wire and_not_n1058_n1061;
    wire not_n1230;
    wire and_not_n379_4_not_n957;
    wire and_not_pi129_138412872010_not_n685;
    wire not_pi048_3;
    wire n562;
    wire n847;
    wire n639;
    wire n1523;
    wire not_pi021_2;
    wire po063_driver;
    wire not_pi003_403536070;
    wire and_pi137_not_n1526;
    wire not_pi051;
    wire not_n988;
    wire not_n544;
    wire and_not_pi009_5_not_pi010_3;
    wire and_not_pi129_103677930763188441902487387275962551382129494864490_not_n1393;
    wire and_not_n1342_not_n1343;
    wire and_pi082_n1582;
    wire n1281;
    wire and_n448_n631;
    wire and_not_pi116_9_n1192;
    wire n1330;
    wire not_n883;
    wire n501;
    wire and_not_n975_n980;
    wire n911;
    wire n578;
    wire n676;
    wire and_not_pi129_10045252112690790399992215344966975021805416861747224664747430_not_n1571;
    wire not_n809;
    wire n1547;
    wire and_pi022_not_pi054_168070;
    wire and_not_n1019_not_n1022;
    wire po011_driver;
    wire and_n390_n403;
    wire not_n1346;
    wire and_not_pi043_2_n387;
    wire not_pi053_1;
    wire not_n540;
    wire not_pi138_6;
    wire n1372;
    wire not_n766;
    wire not_pi021_3;
    wire and_not_pi129_273687473400809163430_not_n894;
    wire and_not_pi027_490_not_n1226;
    wire not_pi054_8235430;
    wire po010_driver;
    wire n1324;
    wire not_n1512;
    wire not_n804;
    wire and_pi064_n1071;
    wire not_pi129_1915812313805664144010;
    wire not_pi026_2;
    wire not_n863;
    wire n655;
    wire and_not_pi039_n722;
    wire not_n718;
    wire and_pi028_not_n798;
    wire and_pi028_n442;
    wire n979;
    wire and_not_pi015_0_n573;
    wire n786;
    wire or_pi129_n1159;
    wire n1265;
    wire n1594;
    wire n350;
    wire and_not_pi027_1_not_pi085_3;
    wire n1147;
    wire and_n1192_n1200;
    wire not_n1080;
    wire and_n301_not_n328;
    wire and_n724_n1146;
    wire and_not_pi027_3_n713;
    wire not_n921;
    wire n1606;
    wire and_not_n718_not_n738;
    wire not_n1423_1;
    wire and_not_pi129_70_not_n541;
    wire not_n1352;
    wire not_n910;
    wire po107_driver;
    wire and_not_pi003_6_n532;
    wire n766;
    wire n1450;
    wire and_not_pi139_n1249;
    wire n1515;
    wire n859;
    wire not_n507;
    wire not_n1287;
    wire and_pi036_n1360;
    wire and_not_pi129_1742514982336908143055105517947102601079450420187483430_not_n1417;
    wire not_n1539;
    wire po045_driver;
    wire and_n927_n1006;
    wire n305;
    wire n1437;
    wire n1175;
    wire and_not_n1205_not_n1208;
    wire and_n379_not_n986;
    wire not_n1546;
    wire not_pi026_6;
    wire n1610;
    wire n1595;
    wire not_pi053_0;
    wire n1489;
    wire and_pi085_pi116;
    wire not_pi026_3430;
    wire and_pi080_not_pi138_3430;
    wire n1500;
    wire and_not_pi129_not_n338;
    wire n990;
    wire n1616;
    wire po098_driver;
    wire not_pi142_0;
    wire n346;
    wire not_pi129_1070069044235980333563563003849377848070;
    wire n1415;
    wire and_not_pi012_n295;
    wire n845;
    wire n836;
    wire and_n379_not_n950;
    wire n974;
    wire and_not_pi005_2_n450;
    wire n680;
    wire n1375;
    wire and_not_n1594_not_n1596;
    wire not_n1049;
    wire and_n934_n1042;
    wire and_n356_n622;
    wire and_not_pi129_405362155971443868320658661090166738008752222510120837461924544480010_not_n1620;
    wire n667;
    wire n1029;
    wire not_pi027_490;
    wire n1555;
    wire and_not_pi129_6782230728490_not_n758;
    wire n1446;
    wire and_not_pi003_5585458640832840070_n1598;
    wire and_n990_n1105;
    wire not_n850;
    wire and_not_n1474_not_n1475;
    wire n1440;
    wire not_pi138_168070;
    wire n359;
    wire and_not_pi007_3_not_n360;
    wire and_pi137_not_n1472;
    wire and_n503_n505;
    wire not_pi013;
    wire not_n1444;
    wire and_not_n379_0_not_n576;
    wire and_not_pi017_4_not_pi018_2;
    wire not_pi050_4;
    wire not_n791;
    wire not_n534;
    wire not_n1507;
    wire n1123;
    wire n1050;
    wire not_n1008;
    wire n1462;
    wire and_pi072_n994;
    wire po043_driver;
    wire n1332;
    wire and_not_pi007_7_n417;
    wire and_n1073_n1075;
    wire not_n1367;
    wire or_pi129_n1298;
    wire and_not_pi129_2569235775210588780886114772242356213216070_not_n1332;
    wire and_n464_n467;
    wire not_n523;
    wire not_n1272;
    wire and_n515_n562;
    wire n975;
    wire not_pi129_2569235775210588780886114772242356213216070;
    wire not_n321;
    wire not_n1372;
    wire and_not_pi110_5_n1369;
    wire n751;
    wire n689;
    wire n1058;
    wire not_n1461;
    wire and_not_pi129_70316764788835532799945507414768825152637918032230572653232010_not_n1576;
    wire not_pi129;
    wire n1231;
    wire and_not_pi063_pi136;
    wire n372;
    wire not_n557;
    wire po099_driver;
    wire and_n1250_n1251;
    wire not_n815;
    wire n1302;
    wire not_n1316;
    wire n861;
    wire n455;
    wire n723;
    wire n894;
    wire and_pi136_pi137;
    wire and_not_n890_not_n891;
    wire not_n794;
    wire and_n638_n990;
    wire and_not_n1222_not_n1225;
    wire and_not_pi096_0_n763;
    wire n735;
    wire and_not_pi129_5_not_n469;
    wire n1475;
    wire and_not_pi003_24010_n670;
    wire and_not_n379_3430_not_n1102;
    wire n1400;
    wire n770;
    wire not_pi003_4;
    wire not_n1508;
    wire not_pi059;
    wire n364;
    wire and_n488_n489;
    wire po004_driver;
    wire n788;
    wire and_not_pi129_403536070_not_n660;
    wire not_n486;
    wire not_n425;
    wire or_pi129_n1263;
    wire not_n729;
    wire n1576;
    wire not_n1348;
    wire not_n949;
    wire n682;
    wire not_pi017_3;
    wire not_n1517;
    wire and_not_n755_not_n843;
    wire and_not_pi008_2_not_pi017_2;
    wire and_not_pi053_6_not_n1173;
    wire and_n503_n559;
    wire and_not_pi129_113988951853731430_not_n866;
    wire not_n1488;
    wire and_not_pi077_not_pi138_5;
    wire and_not_pi011_6_not_pi022_4;
    wire and_not_pi129_4599865365447399609768010_not_n945;
    wire n1293;
    wire n491;
    wire n1556;
    wire n356;
    wire and_not_n713_0_not_n1530;
    wire not_n1082;
    wire n818;
    wire and_not_pi065_0_not_pi138_6;
    wire not_n1407;
    wire n677;
    wire not_n1534;
    wire n329;
    wire and_n379_not_n1082;
    wire not_n1325_3;
    wire n1452;
    wire and_not_n1500_not_n1501;
    wire n408;
    wire n1105;
    wire n1146;
    wire not_pi129_168830552257994114252669163302859949191483641195385604940410056010;
    wire not_n1516;
    wire n1148;
    wire and_n390_n706;
    wire not_n1518;
    wire n1399;
    wire not_pi129_26517308458596534717790233816010;
    wire not_n783;
    wire n358;
    wire po134_driver;
    wire not_pi024_0;
    wire not_n1544;
    wire n791;
    wire n1428;
    wire and_not_pi012_2_n461;
    wire n1261;
    wire and_n638_n642;
    wire n744;
    wire not_n816;
    wire not_pi129_1299348114471230201171721456984490;
    wire not_n1451;
    wire n785;
    wire and_not_pi056_0_not_n301;
    wire not_n511;
    wire n1429;
    wire not_n1339;
    wire and_not_n805_not_n806;
    wire not_n414;
    wire and_pi014_not_pi054_9;
    wire not_n1490;
    wire not_n1067;
    wire not_pi040;
    wire n1140;
    wire and_not_n933_n937;
    wire and_pi011_not_pi054_6;
    wire not_pi054_24010;
    wire and_not_n1053_n1062;
    wire n1009;
    wire and_not_n1231_not_n1232;
    wire not_pi129_492217353521848729599618551903381776068465426225614008572624070;
    wire n330;
    wire not_pi026_1;
    wire and_n503_n513;
    wire not_pi106_4;
    wire not_pi106_0;
    wire not_pi006;
    wire and_n934_n935;
    wire po057_driver;
    wire not_n1524;
    wire not_pi116_5;
    wire and_not_pi003_332329305696010_n1373;
    wire and_n389_n1012;
    wire not_n1050;
    wire and_not_pi096_3_n1145;
    wire n1522;
    wire and_n479_n678;
    wire n523;
    wire n832;
    wire not_n1301;
    wire and_not_pi058_3_not_n835;
    wire and_n347_n417;
    wire not_pi116_0;
    wire n434;
    wire not_pi129_43181145673964365640352930977077280875522488490;
    wire n608;
    wire not_pi019;
    wire and_pi092_pi138;
    wire n1477;
    wire not_n720;
    wire not_n836;
    wire or_n1457_n1464;
    wire not_n940;
    wire and_not_pi013_5_n450;
    wire and_not_pi025_0_pi029;
    wire not_pi044_3;
    wire not_n1502;
    wire and_n446_n453;
    wire n472;
    wire n1476;
    wire and_not_n379_70_not_n1070;
    wire n1159;
    wire not_n1166;
    wire n644;
    wire not_n1020;
    wire not_pi136_10;
    wire n858;
    wire and_not_pi129_332329305696010_not_n784;
    wire n955;
    wire n302;
    wire po032_driver;
    wire not_pi022_1;
    wire n480;
    wire not_pi129_11044276742439206463052992010;
    wire and_not_n897_not_n898;
    wire not_n1433;
    wire n1101;
    wire and_not_n1545_not_n1546;
    wire n342;
    wire n558;
    wire not_n1276;
    wire and_not_pi038_not_pi050;
    wire not_n797;
    wire not_n1423_2;
    wire po097_driver;
    wire n1091;
    wire po088_driver;
    wire not_pi129_0;
    wire n548;
    wire not_n578;
    wire n1527;
    wire not_n865;
    wire not_n1168;
    wire and_not_pi010_1_n449;
    wire not_pi138_10;
    wire and_pi026_n855;
    wire or_pi003_not_n339;
    wire and_not_pi095_not_pi100;
    wire not_n965;
    wire n1015;
    wire and_not_n357_not_n358;
    wire n423;
    wire and_n611_n614;
    wire not_n1563;
    wire not_pi058_10;
    wire not_n658;
    wire and_pi082_not_n1030;
    wire not_pi070;
    wire not_pi073;
    wire not_pi007_4;
    wire and_n408_n1001;
    wire not_n1392;
    wire n875;
    wire n717;
    wire not_n1167;
    wire n1583;
    wire and_n487_n493;
    wire and_pi054_n300;
    wire and_not_n1420_not_n1422;
    wire and_pi025_not_pi116;
    wire n1426;
    wire and_not_n947_not_n951;
    wire and_n737_n1207;
    wire not_n1590;
    wire not_n520;
    wire not_n1347;
    wire n1497;
    wire not_n468;
    wire not_n365;
    wire and_n774_n1374;
    wire not_n1335;
    wire and_not_pi047_1_n568;
    wire not_pi137_70;
    wire and_n579_n919;
    wire n1280;
    wire not_n835;
    wire and_not_n672_not_n681;
    wire not_pi003_9;
    wire n581;
    wire n708;
    wire po072_driver;
    wire n1142;
    wire n1225;
    wire po085_driver;
    wire n647;
    wire not_pi129_3445521474652941107197329863323672432479257983579298060008368490;
    wire not_pi129_1742514982336908143055105517947102601079450420187483430;
    wire n910;
    wire and_pi082_not_n390;
    wire not_n646;
    wire not_n1454;
    wire and_not_pi003_8_n555;
    wire n462;
    wire and_not_pi106_not_n863;
    wire not_n779;
    wire and_pi068_not_n1247_3;
    wire not_n1247_1;
    wire not_n1065;
    wire n392;
    wire not_pi116_1;
    wire and_n447_n466;
    wire and_pi058_pi116;
    wire and_not_pi003_968890104070_n1203;
    wire not_n1557;
    wire and_pi137_not_n1549;
    wire n965;
    wire n1300;
    wire and_pi091_not_n1386_2;
    wire and_not_n379_10_not_n1056;
    wire not_n1584;
    wire not_n379_5;
    wire not_pi138_4;
    wire n1479;
    wire and_not_pi136_168070_not_n1547;
    wire and_not_pi053_3_not_n816;
    wire and_n379_not_n693;
    wire n976;
    wire not_pi129_1435036016098684342856030763566710717400773837392460666392490;
    wire po055_driver;
    wire po049_driver;
    wire n1525;
    wire n486;
    wire and_pi007_not_pi054_2;
    wire and_pi088_pi106;
    wire not_n1362;
    wire n1351;
    wire n1316;
    wire n1600;
    wire n1192;
    wire not_n1208;
    wire and_not_n544_not_n553;
    wire and_pi097_n1149;
    wire and_n726_n787;
    wire not_n1222;
    wire and_not_pi002_n391;
    wire not_n1386_3;
    wire n993;
    wire n1509;
    wire and_not_pi045_4_not_n1033;
    wire and_not_n753_not_n757;
    wire n977;
    wire and_n1251_n1270;
    wire not_pi129_185621159210175743024531636712070;
    wire and_not_pi071_0_not_pi138_24010;
    wire po047_driver;
    wire not_n1421;
    wire and_not_n794_0_not_n1570;
    wire n824;
    wire and_pi143_n1414;
    wire not_n1620;
    wire n1313;
    wire and_pi043_n641;
    wire n1539;
    wire not_pi012_5;
    wire n802;
    wire not_pi137_1;
    wire not_n822;
    wire and_n416_n527;
    wire and_pi059_not_pi116_70;
    wire n487;
    wire n1620;
    wire n1256;
    wire and_pi090_not_n1386_1;
    wire and_not_pi005_not_pi022;
    wire n933;
    wire not_pi106;
    wire n1629;
    wire and_not_n498_not_n507;
    wire and_n398_n401;
    wire and_not_pi129_4_not_n455;
    wire and_not_pi003_2_n484;
    wire not_pi058_1;
    wire n631;
    wire and_pi082_not_pi137_3;
    wire n882;
    wire n313;
    wire and_not_pi012_5_n606;
    wire po066_driver;
    wire not_n1331;
    wire and_n344_n561;
    wire and_not_pi017_not_pi021;
    wire n1233;
    wire not_n1343;
    wire and_not_n1040_n1045;
    wire and_pi122_pi127;
    wire and_n526_n529;
    wire and_pi028_not_pi116_3;
    wire not_n1152;
    wire n725;
    wire not_n1125;
    wire not_pi140_0;
    wire not_n1442;
    wire and_pi094_not_n1167;
    wire n1490;
    wire n431;
    wire not_n1068;
    wire po015_driver;
    wire not_pi011_4;
    wire and_not_pi024_1_n380;
    wire not_n725;
    wire n1210;
    wire po060_driver;
    wire and_not_pi003_47475615099430_n1234;
    wire and_pi006_not_pi054_1;
    wire not_n1198;
    wire n1170;
    wire n296;
    wire not_pi085_7;
    wire and_not_n657_not_n658;
    wire n804;
    wire n978;
    wire not_pi006_0;
    wire not_n1271_1;
    wire n306;
    wire po050_driver;
    wire not_n553;
    wire not_pi053_3;
    wire not_pi053_7;
    wire n843;
    wire not_pi068;
    wire and_not_pi129_3119734822845423713013303218219760490_not_n1152;
    wire and_pi100_pi138;
    wire not_n1386_0;
    wire po065_driver;
    wire and_pi089_not_n1386_0;
    wire and_not_n1473_not_n1477;
    wire and_pi063_n702;
    wire not_n896;
    wire not_n961;
    wire and_not_pi136_57648010_pi139;
    wire not_n952;
    wire and_pi111_not_n1421_0;
    wire po048_driver;
    wire not_pi038_0;
    wire po071_driver;
    wire not_n846;
    wire and_pi033_not_pi109_2;
    wire and_n609_n615;
    wire n433;
    wire n1305;
    wire and_not_n726_0_not_n792;
    wire and_pi041_pi082;
    wire and_n838_n843;
    wire not_n1010;
    wire not_n1022;
    wire and_n390_n960;
    wire not_n334;
    wire and_not_pi038_2_n641;
    wire not_pi129_21838143759917965991093122527538323430;
    wire or_n1237_n1238;
    wire not_pi129_490;
    wire and_pi069_not_n1247_4;
    wire and_pi077_not_n1271_6;
    wire and_not_pi144_0_n1271;
    wire not_pi129_29286449308136415160327158440136953416342323212091034008010;
    wire n1531;
    wire not_pi129_63668057609090279857414351392240010;
    wire and_not_n1272_not_n1273;
    wire not_n1170;
    wire po118_driver;
    wire n1219;
    wire po023_driver;
    wire n1485;
    wire not_pi054_5;
    wire n353;
    wire not_n1463;
    wire n985;
    wire not_n945;
    wire not_pi129_2115876138024253916377293617876786762900601936010;
    wire not_n849;
    wire not_pi129_17984650426474121466202803405696493492512490;
    wire and_pi000_not_pi123;
    wire n535;
    wire n525;
    wire n1361;
    wire not_pi013_3;
    wire not_n1109;
    wire not_pi106_9;
    wire not_n1325_5;
    wire and_n499_n501;
    wire not_n1553;
    wire and_not_pi009_2_n449;
    wire and_not_pi024_3_n692;
    wire n864;
    wire n1512;
    wire not_pi054_490;
    wire not_n695;
    wire and_not_n595_not_n600;
    wire and_pi119_pi138;
    wire n1049;
    wire n1628;
    wire and_not_pi011_4_n418;
    wire n816;
    wire and_not_pi129_1299348114471230201171721456984490_not_n1117;
    wire not_n913;
    wire n1129;
    wire n1516;
    wire not_n1613;
    wire n335;
    wire not_n458;
    wire not_n1325;
    wire and_pi076_not_n1271_5;
    wire not_pi022_3;
    wire and_pi057_not_pi058_9;
    wire and_pi027_pi116;
    wire and_not_pi027_8_pi028;
    wire n731;
    wire n416;
    wire n737;
    wire n1255;
    wire not_pi129_5;
    wire and_not_n379_490_not_n1090;
    wire not_pi129_5080218607396233653221881976522165017724345248360010;
    wire and_not_pi006_not_pi007;
    wire and_not_pi009_4_pi013;
    wire not_n893;
    wire n1352;
    wire and_not_n1114_not_n1115;
    wire not_pi029;
    wire and_not_pi129_21838143759917965991093122527538323430_not_n1184;
    wire n484;
    wire not_pi077;
    wire n899;
    wire not_pi138_1176490;
    wire po068_driver;
    wire not_pi023;
    wire n970;
    wire not_pi137_4;
    wire n1535;
    wire n1187;
    wire not_n307;
    wire not_n1597;
    wire not_pi085_3;
    wire and_pi050_n1041;
    wire n1321;
    wire po106_driver;
    wire not_n483;
    wire and_not_pi003_168070_n683;
    wire not_n825;
    wire and_not_pi129_43181145673964365640352930977077280875522488490_not_n1372;
    wire not_n1247;
    wire not_n1434;
    wire n706;
    wire po028_driver;
    wire n1117;
    wire n311;
    wire not_pi008_0;
    wire and_n379_not_n921;
    wire not_n1500;
    wire and_not_pi003_2326305139872070_not_n1246;
    wire and_not_pi026_4_not_n723_0;
    wire not_n951;
    wire not_n1066;
    wire not_n1382;
    wire not_pi145;
    wire not_n1112;
    wire not_n1409;
    wire not_pi076;
    wire not_pi136_3;
    wire n917;
    wire not_pi129_14811132966169777414641055325137507340304213552070;
    wire not_pi024_4;
    wire and_not_pi129_302268019717750559482470516839540966128657419430_not_n1379;
    wire and_not_pi017_0_n330;
    wire not_pi129_7490483309651862334944941026945644936490;
    wire n400;
    wire and_not_pi026_8_n749;
    wire and_n418_n422;
    wire not_n700;
    wire n1122;
    wire not_n1189;
    wire not_n1101;
    wire and_n772_n774;
    wire and_pi049_not_n1107;
    wire n355;
    wire not_n360;
    wire n399;
    wire n1087;
    wire n1359;
    wire n584;
    wire n808;
    wire not_n1305;
    wire not_pi129_3788186922656647816827176259430;
    wire and_not_pi027_9_not_n845;
    wire not_n1031;
    wire and_n302_not_n334;
    wire and_not_n903_not_n907;
    wire not_n1330;
    wire and_pi018_n295;
    wire not_pi129_39098210485829880490;
    wire n596;
    wire and_pi037_not_pi116_8;
    wire n1529;
    wire n871;
    wire n534;
    wire n1578;
    wire n762;
    wire not_pi047_2;
    wire not_pi116_6;
    wire n662;
    wire not_n904;
    wire not_n1387;
    wire not_n371;
    wire and_not_pi053_not_n745;
    wire n750;
    wire not_pi003_490;
    wire and_pi120_pi138;
    wire and_not_pi003_273687473400809163430_n1619;
    wire not_n1445;
    wire and_not_pi064_not_pi138_8235430;
    wire not_n1142;
    wire and_pi139_n1386;
    wire n1317;
    wire not_n817;
    wire n913;
    wire and_pi082_not_n1028;
    wire and_pi035_pi109;
    wire and_not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070_n1623;
    wire not_n1416;
    wire po036_driver;
    wire and_pi058_not_n839;
    wire n1113;
    wire not_pi006_3;
    wire not_n957;
    wire not_n966;
    wire and_not_pi050_4_not_n1124;
    wire n690;
    wire and_not_pi096_4_pi125;
    wire and_pi016_pi054;
    wire po124_driver;
    wire n1374;
    wire not_n1422;
    wire n473;
    wire not_n408;
    wire not_pi137_5;
    wire n705;
    wire not_n1277;
    wire and_pi034_pi136;
    wire and_not_pi138_9_not_n1493;
    wire not_n1576;
    wire not_pi129_19773267430;
    wire n1011;
    wire not_n1236;
    wire po031_driver;
    wire and_pi018_not_pi054_490;
    wire n1249;
    wire and_not_n1552_not_n1553;
    wire n715;
    wire n563;
    wire n914;
    wire and_n478_n481;
    wire not_n1033;
    wire and_n1246_not_n1591;
    wire and_not_pi129_57648010_not_n635;
    wire not_pi054_4;
    wire n793;
    wire not_n1428;
    wire and_not_pi129_9095436801298611408202050198891430_not_n1132;
    wire and_pi116_not_n796_0;
    wire and_not_n1191_not_n1193;
    wire not_pi071_0;
    wire and_pi062_not_n1247;
    wire n1102;
    wire n385;
    wire and_not_n989_n998;
    wire n1588;
    wire and_pi096_not_n1423_0;
    wire n511;
    wire n1196;
    wire and_not_pi050_1_n403;
    wire po140_driver;
    wire and_pi005_not_pi007_9;
    wire not_pi050_0;
    wire n749;
    wire and_not_n1444_not_n1445;
    wire n1054;
    wire n820;
    wire n848;
    wire and_n386_n393;
    wire and_pi082_not_n948;
    wire not_n1477;
    wire and_pi138_not_n1468;
    wire and_pi084_not_pi136_70;
    wire and_n1100_not_n1109;
    wire n921;
    wire not_n379_168070;
    wire n1287;
    wire and_not_n1377_not_n1378;
    wire not_pi065;
    wire and_not_n1125_n1134;
    wire and_not_n379_1_not_n646;
    wire and_not_n1562_not_n1563;
    wire n1466;
    wire n580;
    wire and_not_po129_n1162;
    wire not_n1218;
    wire not_n1571;
    wire and_n345_n597;
    wire not_pi038_2;
    wire po135_driver;
    wire not_pi142;
    wire not_pi110_1;
    wire n928;
    wire not_n1309;
    wire not_n1537;
    wire and_pi141_n1386;
    wire not_n541;
    wire and_n445_n608;
    wire and_not_n904_not_n905;
    wire n1108;
    wire and_n942_not_n944;
    wire and_n345_n357;
    wire n898;
    wire and_not_pi026_3_n787;
    wire and_not_n310_not_n333;
    wire and_not_pi136_24010_not_n1540;
    wire not_pi026_3;
    wire n900;
    wire and_not_n314_not_n315;
    wire and_pi020_n411;
    wire not_pi085_10;
    wire and_not_pi049_0_n383;
    wire n1240;
    wire n1309;
    wire not_n1504;
    wire not_pi061;
    wire and_pi082_not_n1049;
    wire n924;
    wire and_pi025_not_pi029_0;
    wire and_n406_n579;
    wire not_n889;
    wire not_n554;
    wire not_n1119;
    wire not_n1069;
    wire n1557;
    wire not_n1547;
    wire n401;
    wire and_n432_n434;
    wire and_pi060_not_n1236;
    wire and_pi054_not_n305;
    wire and_n612_n613;
    wire and_n450_n621;
    wire and_not_n313_not_n319;
    wire and_n299_n665;
    wire n572;
    wire and_not_pi009_not_pi011;
    wire and_not_pi039_0_not_pi052_0;
    wire and_not_pi058_0_n773;
    wire not_n831;
    wire n1164;
    wire not_n682;
    wire and_n300_not_n371;
    wire n842;
    wire and_not_pi106_7_not_n941;
    wire n496;
    wire and_n399_n704;
    wire n1216;
    wire not_pi012;
    wire and_not_pi038_1_not_n923;
    wire n1051;
    wire po101_driver;
    wire po096_driver;
    wire not_n1608;
    wire not_pi129_2326305139872070;
    wire n1006;
    wire not_pi027_5;
    wire n904;
    wire po089_driver;
    wire n634;
    wire and_n388_n391;
    wire and_not_n1524_not_n1525;
    wire n1157;
    wire not_pi138_5;
    wire and_not_n1130_n1133;
    wire and_not_pi106_2_not_n885;
    wire and_pi015_not_n581;
    wire n1226;
    wire and_not_pi146_n1249;
    wire n1183;
    wire not_n1491;
    wire n740;
    wire and_not_pi113_n426;
    wire not_n1313;
    wire and_not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430_not_n1629;
    wire not_pi058_3;
    wire and_n934_n1011;
    wire n557;
    wire n826;
    wire not_n1567;
    wire and_not_pi142_0_n1271;
    wire n611;
    wire n1012;
    wire and_not_n307_not_n337;
    wire and_not_n1451_not_n1455;
    wire and_not_pi069_0_pi136;
    wire not_pi012_1;
    wire and_not_pi003_403536070_n827;
    wire n1014;
    wire and_not_n397_not_n413;
    wire n599;
    wire not_n324;
    wire and_pi036_not_pi109_5;
    wire and_n459_n462;
    wire and_not_n1589_not_n1590;
    wire and_pi133_n1631;
    wire and_pi082_not_n972;
    wire not_pi137_7;
    wire n1045;
    wire n673;
    wire not_n887;
    wire not_pi024;
    wire and_not_n728_0_n762;
    wire and_pi095_not_pi096_1;
    wire and_pi081_not_n1325_2;
    wire n1346;
    wire not_n1448;
    wire and_pi005_not_pi054_0;
    wire not_n379_7;
    wire and_pi068_n1039;
    wire po022_driver;
    wire n1154;
    wire and_n416_n430;
    wire n686;
    wire not_n352;
    wire and_not_n1521_not_n1522;
    wire and_pi015_n411;
    wire and_not_n1440_not_n1441;
    wire n931;
    wire and_not_n761_0_not_n1371;
    wire and_not_pi136_2_not_n1358;
    wire not_n1440;
    wire not_pi046;
    wire n1291;
    wire n1391;
    wire and_pi139_n1325;
    wire and_pi082_not_n1157;
    wire and_not_pi046_2_not_n1052;
    wire n589;
    wire and_not_pi019_1_n630;
    wire not_n1458;
    wire and_not_pi129_1181813865805958799768684143120019644340385488367699234582870392070_not_n1608;
    wire not_pi046_0;
    wire n398;
    wire and_n301_not_n302;
    wire n716;
    wire and_pi085_not_n812;
    wire not_n620;
    wire and_not_pi129_657123623635342801395430_not_n936;
    wire n1404;
    wire and_not_n410_not_n411;
    wire not_n839;
    wire not_pi129_597682638941559493067901192655856192170251494124306816490;
    wire n412;
    wire not_pi139_0;
    wire n1519;
    wire not_n519;
    wire not_n1255;
    wire not_n1526;
    wire and_not_n590_not_n591;
    wire not_n323;
    wire and_not_pi013_0_not_n317;
    wire not_n654;
    wire and_n1223_n1228;
    wire not_pi129_4183778472590916451475308348590993345191760458870147715430;
    wire and_pi025_not_pi026_1;
    wire not_n375;
    wire and_not_n1092_n1097;
    wire n1623;
    wire n561;
    wire and_pi091_pi106;
    wire not_n1585;
    wire not_n864;
    wire n1040;
    wire not_pi003_70;
    wire not_pi129_16284135979104490;
    wire n1366;
    wire not_n868;
    wire and_n475_n477;
    wire not_pi129_9095436801298611408202050198891430;
    wire or_pi129_n1293;
    wire n730;
    wire n478;
    wire not_n995;
    wire not_pi042;
    wire not_n1386_2;
    wire and_not_pi002_5_n383;
    wire and_not_pi114_pi123;
    wire n792;
    wire n906;
    wire not_n1468;
    wire and_not_pi138_10_not_n1508;
    wire not_n838;
    wire n595;
    wire and_not_n1537_not_n1541;
    wire n307;
    wire not_n1179;
    wire not_n1489;
    wire not_n379_2;
    wire not_pi129_403536070;
    wire not_pi001;
    wire and_not_pi006_3_n341;
    wire n1542;
    wire not_n1209;
    wire not_n564;
    wire n721;
    wire n1288;
    wire n1263;
    wire and_pi085_not_pi116_1;
    wire not_n1601;
    wire and_not_pi021_1_n300;
    wire po123_driver;
    wire not_pi141;
    wire and_not_n1403_not_n1404;
    wire not_pi042_2;
    wire and_pi017_n612;
    wire and_not_pi069_n1103;
    wire and_not_n379_24010_not_n1128;
    wire not_pi064;
    wire not_n616;
    wire and_not_pi026_10_n1155;
    wire and_n387_n388;
    wire n795;
    wire and_not_pi116_4_n818;
    wire and_pi019_n664;
    wire po038_driver;
    wire not_pi010;
    wire and_n298_n299;
    wire and_not_n861_not_n862;
    wire not_pi044_1;
    wire and_not_pi009_0_not_n367;
    wire n1421;
    wire and_pi030_n1360;
    wire n1503;
    wire and_n448_n465;
    wire and_not_pi129_492217353521848729599618551903381776068465426225614008572624070_n1586;
    wire and_not_pi016_1_n354;
    wire not_pi046_2;
    wire and_n503_n674;
    wire and_n649_n707;
    wire not_n1381;
    wire not_n713_0;
    wire n587;
    wire not_n379_3;
    wire and_pi052_not_n940_0;
    wire and_pi132_pi133;
    wire and_not_pi129_125892552985318850263419623839875454447587430_not_n1340;
    wire and_pi090_n1249;
    wire and_n447_n452;
    wire and_n724_not_n833;
    wire not_pi136_6;
    wire and_not_n1168_not_n1172;
    wire n641;
    wire n1526;
    wire and_not_pi029_1_pi059;
    wire not_pi028_1;
    wire not_pi065_0;
    wire not_n1496;
    wire not_n435;
    wire n1195;
    wire not_pi048;
    wire n1363;
    wire n813;
    wire and_not_n1387_not_n1388;
    wire and_not_n379_7_not_n1008;
    wire and_not_pi137_4_not_n1456;
    wire and_n514_n518;
    wire and_not_n1304_not_n1305;
    wire and_n459_n479;
    wire not_n1151;
    wire and_pi073_not_n1271_2;
    wire not_n350;
    wire and_not_n1365_not_n1366;
    wire not_n956;
    wire not_n1193;
    wire and_n638_n1027;
    wire and_not_n1346_not_n1347;
    wire not_pi053_8;
    wire n1548;
    wire and_pi082_not_n700;
    wire and_pi136_not_n1554;
    wire n1448;
    wire not_pi129_332329305696010;
    wire n1532;
    wire n1621;
    wire not_n1205;
    wire not_pi009_3;
    wire not_pi106_7;
    wire and_n389_n392;
    wire not_n1028;
    wire and_not_n842_not_n844;
    wire n709;
    wire and_pi027_n838;
    wire po131_driver;
    wire n886;
    wire n1232;
    wire and_not_pi048_1_n381;
    wire and_not_n379_3_not_n931;
    wire not_n767;
    wire po132_driver;
    wire and_pi060_n1144;
    wire and_not_pi026_7_not_pi027_7;
    wire and_not_pi005_3_not_pi007_5;
    wire not_pi017_0;
    wire not_pi041_2;
    wire and_pi082_not_n1037;
    wire not_n305;
    wire n1077;
    wire and_n356_n433;
    wire not_n325;
    wire not_n366;
    wire and_n400_n401;
    wire n437;
    wire n1130;
    wire and_n1251_n1261;
    wire n1534;
    wire not_n1628;
    wire po069_driver;
    wire n1013;
    wire po017_driver;
    wire n1546;
    wire not_pi058_8;
    wire n1308;
    wire not_pi022_0;
    wire not_n744;
    wire and_pi100_not_n1423_2;
    wire po130_driver;
    wire and_not_pi014_0_not_n320;
    wire not_n1325_6;
    wire n872;
    wire not_n784;
    wire n600;
    wire and_not_pi129_93874803376477543056490_not_n915;
    wire not_pi027_6;
    wire not_pi003_113988951853731430;
    wire not_n1575;
    wire not_n691;
    wire not_n936;
    wire not_pi002_5;
    wire not_n944;
    wire not_n1199;
    wire n529;
    wire not_pi054_1;
    wire and_n487_n633;
    wire n803;
    wire n524;
    wire not_n854;
    wire not_n672;
    wire po116_driver;
    wire and_not_n917_not_n922;
    wire not_pi143;
    wire not_n877;
    wire and_pi144_n1414;
    wire not_n1312;
    wire not_pi003_10;
    wire not_n790;
    wire and_pi010_not_pi022_1;
    wire n300;
    wire and_n449_n558;
    wire and_n300_n329;
    wire and_not_pi013_4_n417;
    wire and_pi051_not_pi109_7;
    wire n1055;
    wire and_pi080_not_n1325_1;
    wire and_not_pi058_not_n752;
    wire and_not_pi015_2_not_pi049_1;
    wire not_n769;
    wire not_n1201;
    wire and_n434_n599;
    wire not_n692;
    wire and_not_n458_not_n468;
    wire po016_driver;
    wire not_n379_1;
    wire n884;
    wire n554;
    wire and_pi039_not_n943;
    wire n547;
    wire n1038;
    wire and_n398_n925;
    wire not_pi138_3;
    wire not_pi136_70;
    wire n972;
    wire not_n734;
    wire n812;
    wire not_n953;
    wire n463;
    wire n1082;
    wire n629;
    wire and_not_pi129_47475615099430_not_n770;
    wire not_pi016;
    wire n1434;
    wire n1162;
    wire not_n1429;
    wire not_pi116_9;
    wire n1178;
    wire not_n1252;
    wire and_not_pi007_1_n311;
    wire n1499;
    wire po067_driver;
    wire and_pi082_not_n1018;
    wire n1563;
    wire not_pi017_4;
    wire not_pi122_0;
    wire and_not_n746_not_n751;
    wire n1100;
    wire and_pi026_n768;
    wire not_pi129_3119734822845423713013303218219760490;
    wire not_pi138_403536070;
    wire and_n787_n1175;
    wire and_pi099_n1249;
    wire not_pi058_2;
    wire and_not_n817_not_n821;
    wire not_n412;
    wire and_not_n802_not_n803;
    wire po125_driver;
    wire not_n1034;
    wire n1405;
    wire n1412;
    wire and_not_pi056_n308;
    wire not_pi003_6;
    wire not_n1535;
    wire n498;
    wire and_not_pi073_not_pi136_10;
    wire n438;
    wire n897;
    wire not_n1386_5;
    wire and_not_pi143_n1271;
    wire n468;
    wire not_pi114;
    wire po105_driver;
    wire not_pi136_4;
    wire n552;
    wire not_n1247_5;
    wire not_pi011_1;
    wire not_n920;
    wire n1007;
    wire n1270;
    wire not_pi137_2;
    wire or_pi129_n1268;
    wire not_n1247_0;
    wire po121_driver;
    wire not_n1393;
    wire not_pi005_1;
    wire po009_driver;
    wire not_pi040_1;
    wire n958;
    wire n1419;
    wire and_not_pi129_205005145156954906122290109080958673914396262484637238056070_not_n1446;
    wire and_not_pi054_8235430_pi118;
    wire n515;
    wire not_pi009_2;
    wire n582;
    wire not_n1357;
    wire and_not_n1466_not_n1467;
    wire n1590;
    wire not_pi003_1915812313805664144010;
    wire n984;
    wire n700;
    wire and_not_pi129_1_not_n414;
    wire and_not_pi129_881247870897231951843937366879128181133112010_not_n1344;
    wire and_not_n723_not_n729;
    wire not_pi025_0;
    wire po008_driver;
    wire and_not_pi007_8_n346;
    wire not_n1326;
    wire and_n447_n546;
    wire n428;
    wire n1295;
    wire and_not_pi137_5_not_n1476;
    wire and_not_pi129_63668057609090279857414351392240010_not_n1138;
    wire not_n872;
    wire and_not_pi129_17984650426474121466202803405696493492512490_not_n1336;
    wire and_pi082_not_n1007;
    wire not_n1399;
    wire not_n1415;
    wire and_not_pi129_5080218607396233653221881976522165017724345248360010_not_n1401;
    wire not_n931;
    wire and_not_n1407_not_n1408;
    wire not_pi015_0;
    wire and_not_pi129_24010_not_n593;
    wire not_pi129_12197604876358357001385738625629718207556152941312384010;
    wire and_not_pi100_0_not_n781;
    wire and_n408_n1036;
    wire po025_driver;
    wire not_n409;
    wire not_n1325_2;
    wire and_pi079_not_pi136_6;
    wire and_not_n309_not_n335;
    wire n448;
    wire not_n588;
    wire not_n811;
    wire and_not_n850_not_n852;
    wire and_pi082_not_n589;
    wire not_pi018_2;
    wire not_n793;
    wire not_pi138_2;
    wire not_pi129_8235430;
    wire n291;
    wire not_n1089;
    wire n1209;
    wire and_not_pi106_5_not_n906;
    wire and_pi040_pi082;
    wire po139_driver;
    wire n1552;
    wire n1252;
    wire and_n445_n463;
    wire not_pi111;
    wire and_not_pi129_35561530251773635572553173835655155124070416738520070_not_n1405;
    wire and_not_pi136_4_not_n1450;
    wire not_pi109_6;
    wire n827;
    wire not_n897;
    wire n451;
    wire not_n1340;
    wire n422;
    wire n1567;
    wire not_pi129_405362155971443868320658661090166738008752222510120837461924544480010;
    wire and_not_pi129_6_not_n483;
    wire not_n989;
    wire n1347;
    wire n1601;
    wire not_n741;
    wire n569;
    wire n947;
    wire and_n1251_n1291;
    wire not_pi096_3;
    wire not_pi050_1;
    wire and_pi031_pi109;
    wire n366;
    wire n420;
    wire and_not_pi129_168830552257994114252669163302859949191483641195385604940410056010_n1604;
    wire n885;
    wire and_pi142_n1386;
    wire not_pi024_3;
    wire not_pi097;
    wire and_not_pi129_7490483309651862334944941026945644936490_not_n1233;
    wire n421;
    wire and_not_pi129_3_not_n437;
    wire and_not_pi045_1_n384;
    wire n592;
    wire n1348;
    wire and_not_pi027_3430_n1529;
    wire n754;
    wire and_not_n1399_not_n1400;
    wire n500;
    wire n1498;
    wire n349;
    wire and_not_pi040_n390;
    wire n643;
    wire po035_driver;
    wire not_pi129_541169560379521116689596608490;
    wire and_n301_n302;
    wire not_n1164_0;
    wire not_pi043_1;
    wire and_n754_n787;
    wire not_pi014_1;
    wire n368;
    wire and_n341_n419;
    wire n674;
    wire n427;
    wire n833;
    wire n1111;
    wire not_pi004;
    wire and_not_n1515_not_n1516;
    wire and_not_pi129_3788186922656647816827176259430_not_n1060;
    wire and_n550_n551;
    wire not_n1007;
    wire and_pi034_pi109;
    wire not_n1060;
    wire n1083;
    wire not_n1177;
    wire not_n911;
    wire n1326;
    wire not_n1438;
    wire and_n448_n524;
    wire not_pi129_657123623635342801395430;
    wire and_not_pi026_5_pi027;
    wire and_not_pi110_1_not_n761;
    wire not_pi027;
    wire n1613;
    wire n388;
    wire not_n1503;
    wire n377;
    wire and_n748_n750;
    wire n1124;
    wire not_n1558;
    wire and_not_pi136_5_not_n1461;
    wire and_not_pi129_248930711762415449007872216849586085868492917169640490_not_n1409;
    wire n1469;
    wire n850;
    wire n1474;
    wire n436;
    wire n688;
    wire not_n726_1;
    wire n1507;
    wire and_not_n727_not_n728;
    wire and_pi017_not_pi054_70;
    wire po092_driver;
    wire not_pi106_8;
    wire n930;
    wire n386;
    wire not_n1147;
    wire and_pi136_not_n1536;
    wire not_pi062;
    wire not_pi106_3;
    wire and_not_n325_not_n327;
    wire n426;
    wire not_pi129_4599865365447399609768010;
    wire n622;
    wire and_not_pi129_541169560379521116689596608490_not_n1044;
    wire po091_driver;
    wire not_n582;
    wire and_not_n794_not_n795;
    wire not_n1271;
    wire not_n1136;
    wire n1032;
    wire and_pi088_pi138;
    wire and_not_pi046_0_not_pi050_0;
    wire and_not_pi024_not_pi049;
    wire n1144;
    wire n363;
    wire n446;
    wire and_not_n628_not_n634;
    wire n796;
    wire n1173;
    wire and_not_pi027_70_not_n1198;
    wire and_not_pi137_10_not_n1560;
    wire not_pi129_85383234134508499009700170379408027452893070589186688070;
    wire and_not_pi026_24010_not_n1230;
    wire not_pi026;
    wire not_n730;
    wire not_n894;
    wire po029_driver;
    wire n1411;
    wire n853;
    wire not_n1083;
    wire and_not_pi070_0_not_pi138_70;
    wire not_pi009_1;
    wire n838;
    wire and_n934_n1131;
    wire and_not_pi112_0_not_n1421_1;
    wire po077_driver;
    wire and_not_pi129_16284135979104490_not_n858;
    wire not_n1171;
    wire not_n1523;
    wire not_n1594;
    wire not_n906;
    wire n1598;
    wire not_pi012_0;
    wire and_not_pi003_138412872010_n1185;
    wire n1377;
    wire n830;
    wire not_pi109_2;
    wire and_not_pi002_3_n399;
    wire and_pi082_not_n1101;
    wire n1458;
    wire and_pi024_pi082;
    wire n944;
    wire not_pi138_7;
    wire and_n583_n704;
    wire n695;
    wire not_pi024_2;
    wire not_n842;
    wire n1401;
    wire n1310;
    wire and_not_pi051_0_n736;
    wire n1203;
    wire n520;
    wire not_pi075;
    wire not_n969;
    wire po075_driver;
    wire and_not_n764_not_n765;
    wire and_not_pi058_5_not_pi110_4;
    wire and_not_pi053_5_not_n1148;
    wire and_pi027_n1182;
    wire not_n1325_0;
    wire n1367;
    wire not_n1128;
    wire not_n1327;
    wire and_n1412_n1413;
    wire and_not_pi005_0_not_pi006_1;
    wire n1492;
    wire n692;
    wire and_not_pi106_0_not_n871;
    wire not_n1247_3;
    wire and_n448_n451;
    wire n403;
    wire not_pi054_7;
    wire not_n924;
    wire not_pi054_168070;
    wire n869;
    wire and_n705_n1106;
    wire and_n331_n332;
    wire not_pi085_5;
    wire n1541;
    wire and_n638_n639;
    wire n1420;
    wire n1545;
    wire and_n448_n673;
    wire n943;
    wire not_n901;
    wire and_not_n910_not_n914;
    wire not_n751;
    wire n1107;
    wire not_n761_0;
    wire and_not_pi018_0_n449;
    wire n470;
    wire n1449;
    wire and_not_pi016_2_n351;
    wire not_pi137;
    wire not_n1421_1;
    wire and_not_n782_not_n783;
    wire and_pi012_not_pi054_7;
    wire n896;
    wire not_n810;
    wire n821;
    wire and_not_pi011_2_pi021;
    wire n348;
    wire and_pi011_n459;
    wire n1034;
    wire and_not_n1164_not_n1166;
    wire not_n1220;
    wire n1373;
    wire and_n300_n303;
    wire and_not_pi027_2_not_pi053_1;
    wire and_n838_n856;
    wire and_not_pi116_6_n843;
    wire and_n1175_n1182;
    wire not_pi003_57648010;
    wire n702;
    wire and_not_n604_not_n616;
    wire and_n291_n344;
    wire n703;
    wire not_pi053_2;
    wire not_pi005_3;
    wire n1417;
    wire not_pi136_5;
    wire n568;
    wire n651;
    wire n341;
    wire not_pi116_2;
    wire n338;
    wire not_n1519;
    wire not_pi058_9;
    wire and_pi009_n369;
    wire n1362;
    wire and_pi098_not_n1386_5;
    wire and_not_pi140_n1249;
    wire n615;
    wire not_pi017;
    wire n1199;
    wire n1251;
    wire n868;
    wire not_n310;
    wire not_pi027_8;
    wire not_pi109_7;
    wire n1520;
    wire n779;
    wire n1382;
    wire not_n368;
    wire n616;
    wire and_pi109_n722;
    wire not_n967;
    wire not_n1304;
    wire n1486;
    wire and_n385_n1035;
    wire not_n1115;
    wire or_n1520_n1527;
    wire and_not_n717_not_n719;
    wire not_pi136_2;
    wire not_pi016_0;
    wire not_pi011;
    wire not_n681;
    wire not_pi112_0;
    wire and_not_n423_n424;
    wire not_n379_490;
    wire n458;
    wire not_pi129_6782230728490;
    wire n1061;
    wire not_n1353;
    wire and_not_pi007_10_not_pi009_6;
    wire po074_driver;
    wire not_pi020_0;
    wire n841;
    wire n724;
    wire and_not_pi047_2_n407;
    wire not_n1180;
    wire not_n590;
    wire and_not_n1504_not_n1505;
    wire n316;
    wire not_pi138;
    wire n477;
    wire not_n693;
    wire and_not_pi026_2_n713;
    wire n1153;
    wire not_pi015_2;
    wire po084_driver;
    wire n1151;
    wire n1128;
    wire and_pi027_not_n739;
    wire not_pi137_0;
    wire n488;
    wire not_pi136_1176490;
    wire and_not_pi023_pi055;
    wire not_n1396;
    wire and_pi099_pi106;
    wire and_pi082_not_n1069;
    wire and_pi098_pi138;
    wire not_pi109_5;
    wire n995;
    wire and_not_pi136_not_pi137_1;
    wire and_n1244_n1246;
    wire not_n1481;
    wire not_n1554;
    wire and_pi054_not_n1595;
    wire and_n388_n390;
    wire not_n735;
    wire not_n1521;
    wire n295;
    wire and_n343_n349;
    wire po078_driver;
    wire n1286;
    wire n1481;
    wire not_n1056;
    wire n1125;
    wire and_not_n1308_not_n1309;
    wire n337;
    wire n856;
    wire n963;
    wire not_n738;
    wire and_not_pi041_1_not_pi043_1;
    wire not_pi007_7;
    wire and_n743_n755;
    wire and_not_n831_not_n832;
    wire not_n1164;
    wire not_pi118;
    wire not_n912;
    wire not_n309;
    wire n1060;
    wire and_not_n889_not_n893;
    wire and_not_n435_not_n436;
    wire n1472;
    wire and_pi094_n1324;
    wire n414;
    wire not_n726;
    wire not_n724;
    wire and_not_n440_not_n454;
    wire and_pi116_n1165;
    wire n1297;
    wire n506;
    wire not_pi137_6;
    wire and_pi009_not_pi054_4;
    wire not_n803;
    wire not_n727;
    wire and_pi123_n1236;
    wire not_pi003_3430;
    wire n532;
    wire po020_driver;
    wire n664;
    wire n546;
	INVX1 g_not_pi085_8 (pi085, not_pi085_8);
	INVX1 g_not_pi096_4 (pi096, not_pi096_4);
	AND2X1 g_and_n788_n1370 (n788, n1370, and_n788_n1370);
	AND2X1 g_and_n379_not_n1002 (n379, not_n1002, and_n379_not_n1002);
	INVX1 g_not_n440 (n440, not_n440);
	AND2X1 g_and_pi007_not_n311 (pi007, not_n311, and_pi007_not_n311);
	AND2X1 g_and_not_pi129_2_not_n428 (not_n428, not_pi129_2, and_not_pi129_2_not_n428);
	BUFX2 g_po120 (po120_driver, po120);
	BUFX2 g_n945 (and_n942_not_n944, n945);
	AND2X1 g_and_n704_n1035 (n1035, n704, and_n704_n1035);
	BUFX2 g_n1247 (and_n1244_n1246, n1247);
	AND2X1 g_and_not_n882_not_n886 (not_n882, not_n886, and_not_n882_not_n886);
	INVX1 g_not_pi054_10 (pi054, not_pi054_10);
	BUFX2 g_n1570 (and_not_n737_n795, n1570);
	AND2X1 g_and_not_n1470_not_n1471 (not_n1471, not_n1470, and_not_n1470_not_n1471);
	BUFX2 g_n1456 (and_not_n1451_not_n1455, n1456);
	BUFX2 g_po073 (po073_driver, po073);
	BUFX2 g_n1227 (and_not_pi027_490_not_n1226, n1227);
	BUFX2 g_n636 (and_not_pi129_57648010_not_n635, n636);
	AND2X1 g_and_pi073_n958 (pi073, n958, and_pi073_n958);
	INVX1 g_not_n1460 (n1460, not_n1460);
	BUFX2 g_po070 (po070_driver, po070);
	BUFX2 g_n303 (and_n301_n302, n303);
	INVX1 g_not_n832 (n832, not_n832);
	INVX1 g_not_n1271_2 (n1271, not_n1271_2);
	BUFX2 g_n351 (and_not_pi017_1_pi054, n351);
	AND2X1 g_and_pi086_not_pi138_403536070 (not_pi138_403536070, pi086, and_pi086_not_pi138_403536070);
	INVX1 g_not_n1472 (n1472, not_n1472);
	INVX1 g_not_pi050 (pi050, not_pi050);
	AND2X1 g_and_pi054_not_n336 (not_n336, pi054, and_pi054_not_n336);
	AND2X1 g_and_not_pi129_10_not_n531 (not_pi129_10, not_n531, and_not_pi129_10_not_n531);
	BUFX2 g_n1104 (and_not_pi069_n1103, n1104);
	AND2X1 g_and_not_pi003_3430_n636 (n636, not_pi003_3430, and_not_pi003_3430_n636);
	BUFX2 g_n718 (and_pi025_not_pi116, n718);
	BUFX2 g_n1473 (and_pi137_not_n1472, n1473);
	AND2X1 g_and_not_n1174_not_n1176 (not_n1176, not_n1174, and_not_n1174_not_n1176);
	BUFX2 g_n879 (and_not_pi106_1_not_n878, n879);
	BUFX2 g_n410 (and_pi082_not_n409, n410);
	BUFX2 g_n697 (and_not_pi002_1_not_pi045_3, n697);
	BUFX2 g_n936 (and_n934_n935, n936);
	AND2X1 g_and_not_pi003_7_n542 (n542, not_pi003_7, and_not_pi003_7_n542);
	BUFX2 g_n379 (and_pi122_pi127, n379);
	AND2X1 g_and_not_n1391_not_n1392 (not_n1392, not_n1391, and_not_n1391_not_n1392);
	INVX1 g_not_n1552 (n1552, not_n1552);
	AND2X1 g_and_n385_n697 (n385, n697, and_n385_n697);
	AND2X1 g_and_n754_n755 (n754, n755, and_n754_n755);
	BUFX2 g_n1207 (and_not_pi058_10_n1206, n1207);
	AND2X1 g_and_not_pi138_0_n1246 (not_pi138_0, n1246, and_not_pi138_0_n1246);
	BUFX2 g_n613 (and_not_pi029_1_pi059, n613);
	AND2X1 g_and_not_n1285_not_n1287 (not_n1285, not_n1287, and_not_n1285_not_n1287);
	AND2X1 g_and_pi072_not_n1271_1 (pi072, not_n1271_1, and_pi072_not_n1271_1);
	AND2X1 g_and_not_n1187_not_n1189 (not_n1189, not_n1187, and_not_n1187_not_n1189);
	BUFX2 g_n1416 (and_pi142_n1414, n1416);
	BUFX2 g_po096 (po096_driver, po096);
	INVX1 g_not_n713 (n713, not_n713);
	INVX1 g_not_n1492 (n1492, not_n1492);
	AND2X1 g_and_not_n1218_not_n1220 (not_n1220, not_n1218, and_not_n1218_not_n1220);
	INVX1 g_not_n1187 (n1187, not_n1187);
	INVX1 g_not_n1195 (n1195, not_n1195);
	BUFX2 g_n1030 (and_not_pi024_3_n692, n1030);
	AND2X1 g_and_n398_n399 (n398, n399, and_n398_n399);
	INVX1 g_not_pi054 (pi054, not_pi054);
	AND2X1 g_and_not_pi111_n1621 (n1621, not_pi111, and_not_pi111_n1621);
	AND2X1 g_and_pi059_not_n1217 (pi059, not_n1217, and_pi059_not_n1217);
	BUFX2 g_po066 (po066_driver, po066);
	AND2X1 g_and_n448_n512 (n512, n448, and_n448_n512);
	BUFX2 g_n880 (and_not_n875_not_n879, n880);
	BUFX2 g_n1145 (and_not_pi058_5_not_pi110_4, n1145);
	INVX1 g_not_n1013 (n1013, not_n1013);
	BUFX2 g_n873 (and_not_n868_not_n872, n873);
	BUFX2 g_n625 (and_not_n620_not_n624, n625);
	INVX1 g_not_pi002_1 (pi002, not_pi002_1);
	INVX1 g_not_pi009_5 (pi009, not_pi009_5);
	BUFX2 g_n650 (and_not_pi015_2_not_pi049_1, n650);
	INVX1 g_not_n617 (n617, not_n617);
	INVX1 g_not_pi026_4 (pi026, not_pi026_4);
	AND2X1 g_and_not_pi013_not_pi014 (not_pi013, not_pi014, and_not_pi013_not_pi014);
	INVX1 g_not_n645 (n645, not_n645);
	BUFX2 g_n1478 (and_not_n1473_not_n1477, n1478);
	BUFX2 g_n1540 (and_not_n1538_not_n1539, n1540);
	AND2X1 g_and_pi032_not_pi109_1 (not_pi109_1, pi032, and_pi032_not_pi109_1);
	BUFX2 g_n839 (and_not_n837_not_n838, n839);
	INVX1 g_not_n1004 (n1004, not_n1004);
	AND2X1 g_and_not_pi137_2_not_n1354 (not_n1354, not_pi137_2, and_not_pi137_2_not_n1354);
	AND2X1 g_and_n762_not_n777 (not_n777, n762, and_n762_not_n777);
	BUFX2 g_po129 (po129_driver, po129);
	INVX1 g_not_n575 (n575, not_n575);
	INVX1 g_not_pi058_7 (pi058, not_pi058_7);
	AND2X1 g_and_pi082_not_n409 (not_n409, pi082, and_pi082_not_n409);
	AND2X1 g_and_pi026_pi053 (pi053, pi026, and_pi026_pi053);
	INVX1 g_not_n1215 (n1215, not_n1215);
	BUFX2 g_n304 (and_n300_n303, n304);
	INVX1 g_not_n357 (n357, not_n357);
	INVX1 g_not_n655 (n655, not_n655);
	AND2X1 g_and_not_pi008_n294 (not_pi008, n294, and_not_pi008_n294);
	AND2X1 g_and_pi092_pi106 (pi106, pi092, and_pi092_pi106);
	INVX1 g_not_n1085 (n1085, not_n1085);
	AND2X1 g_and_not_pi008_3_n449 (n449, not_pi008_3, and_not_pi008_3_n449);
	BUFX2 g_n929 (and_n638_n928, n929);
	INVX1 g_not_pi129_152867006319425761937651857692768264010 (pi129, not_pi129_152867006319425761937651857692768264010);
	BUFX2 g_n1245 (and_pi132_pi133, n1245);
	AND2X1 g_and_pi075_not_n1271_4 (not_n1271_4, pi075, and_pi075_not_n1271_4);
	INVX1 g_not_n1497 (n1497, not_n1497);
	AND2X1 g_and_pi116_n1578 (n1578, pi116, and_pi116_n1578);
	INVX1 g_not_n1589 (n1589, not_n1589);
	AND2X1 g_and_not_pi129_725745515342319093317411710931737859674906464051430_not_n1397 (not_pi129_725745515342319093317411710931737859674906464051430, not_n1397, and_not_pi129_725745515342319093317411710931737859674906464051430_not_n1397);
	INVX1 g_not_pi010_3 (pi010, not_pi010_3);
	AND2X1 g_and_pi144_n1386 (n1386, pi144, and_pi144_n1386);
	AND2X1 g_and_not_pi041_0_n405 (n405, not_pi041_0, and_not_pi041_0_n405);
	INVX1 g_not_n332 (n332, not_n332);
	INVX1 g_not_n837 (n837, not_n837);
	AND2X1 g_and_not_n875_not_n879 (not_n875, not_n879, and_not_n875_not_n879);
	AND2X1 g_and_n705_n1100 (n705, n1100, and_n705_n1100);
	AND2X1 g_and_pi095_n1324 (pi095, n1324, and_pi095_n1324);
	BUFX2 g_po126 (po126_driver, po126);
	INVX1 g_not_n1453 (n1453, not_n1453);
	BUFX2 g_n373 (and_n356_n372, n373);
	BUFX2 g_n362 (and_n359_n361, n362);
	INVX1 g_not_pi139 (pi139, not_pi139);
	INVX1 g_not_n907 (n907, not_n907);
	INVX1 g_not_n899 (n899, not_n899);
	INVX1 g_not_n1400 (n1400, not_n1400);
	BUFX2 g_n656 (and_not_n654_not_n655, n656);
	BUFX2 g_n1470 (and_pi079_not_pi136_6, n1470);
	AND2X1 g_and_pi057_not_n1194 (pi057, not_n1194, and_pi057_not_n1194);
	AND2X1 g_and_not_pi129_2824752490_not_n669 (not_n669, not_pi129_2824752490, and_not_pi129_2824752490_not_n669);
	INVX1 g_not_n1379 (n1379, not_n1379);
	BUFX2 g_n1389 (and_not_n1387_not_n1388, n1389);
	INVX1 g_not_pi136_24010 (pi136, not_pi136_24010);
	BUFX2 g_po003 (po003_driver, po003);
	INVX1 g_not_pi044 (pi044, not_pi044);
	INVX1 g_not_n1505 (n1505, not_n1505);
	INVX1 g_not_n1420 (n1420, not_n1420);
	AND2X1 g_and_pi093_pi106 (pi093, pi106, and_pi093_pi106);
	BUFX2 g_n952 (and_not_n947_not_n951, n952);
	BUFX2 g_n1138 (and_not_pi106_8_n1137, n1138);
	BUFX2 g_n1414 (and_n1412_n1413, n1414);
	AND2X1 g_and_n777_n790 (n790, n777, and_n777_n790);
	INVX1 g_not_n870 (n870, not_n870);
	AND2X1 g_and_pi067_not_n1271_0 (pi067, not_n1271_0, and_pi067_not_n1271_0);
	AND2X1 g_and_not_pi015_1_not_n584 (not_pi015_1, not_n584, and_not_pi015_1_not_n584);
	INVX1 g_not_n1538 (n1538, not_n1538);
	INVX1 g_not_pi007_0 (pi007, not_pi007_0);
	INVX1 g_not_n892 (n892, not_n892);
	INVX1 g_not_n1150 (n1150, not_n1150);
	BUFX2 g_n343 (and_n300_n342, n343);
	INVX1 g_not_n379_9 (n379, not_n379_9);
	INVX1 g_not_n624 (n624, not_n624);
	INVX1 g_not_n1113 (n1113, not_n1113);
	INVX1 g_not_pi013_2 (pi013, not_pi013_2);
	BUFX2 g_n800 (and_not_pi026_6_not_pi100_1, n800);
	BUFX2 g_n748 (and_not_pi116_0_n747, n748);
	AND2X1 g_and_n420_n421 (n421, n420, and_n420_n421);
	INVX1 g_not_n1514 (n1514, not_n1514);
	AND2X1 g_and_pi071_not_n1247_6 (pi071, not_n1247_6, and_pi071_not_n1247_6);
	BUFX2 g_po040 (po040_driver, po040);
	AND2X1 g_and_not_n654_not_n655 (not_n654, not_n655, and_not_n654_not_n655);
	AND2X1 g_and_not_n1227_not_n1229 (not_n1229, not_n1227, and_not_n1227_not_n1229);
	INVX1 g_not_n709 (n709, not_n709);
	BUFX2 g_n384 (and_not_pi024_not_pi049, n384);
	BUFX2 g_po114_driver (and_not_pi129_29286449308136415160327158440136953416342323212091034008010_not_n1442, po114_driver);
	INVX1 g_not_n866 (n866, not_n866);
	AND2X1 g_and_not_n965_not_n967 (not_n967, not_n965, and_not_n965_not_n967);
	AND2X1 g_and_n705_n708 (n708, n705, and_n705_n708);
	INVX1 g_not_n1271_6 (n1271, not_n1271_6);
	INVX1 g_not_pi056 (pi056, not_pi056);
	BUFX2 g_po117_driver (or_n1469_n1479, po117_driver);
	BUFX2 g_n1095 (and_n934_n1094, n1095);
	AND2X1 g_and_n445_n480 (n445, n480, and_n445_n480);
	INVX1 g_not_pi096_1 (pi096, not_pi096_1);
	INVX1 g_not_pi021_0 (pi021, not_pi021_0);
	BUFX2 g_po131 (po131_driver, po131);
	BUFX2 g_n513 (and_n448_n512, n513);
	BUFX2 g_n732 (and_not_n730_not_n731, n732);
	BUFX2 g_n811 (and_not_pi100_2_pi116, n811);
	AND2X1 g_and_pi136_not_n1513 (not_n1513, pi136, and_pi136_not_n1513);
	BUFX2 g_n1340 (and_not_n1338_not_n1339, n1340);
	BUFX2 g_po140 (po140_driver, po140);
	AND2X1 g_and_n401_n698 (n698, n401, and_n401_n698);
	INVX1 g_not_n379_6 (n379, not_n379_6);
	OR2X1 g_or_pi129_n1302 (pi129, n1302, or_pi129_n1302);
	INVX1 g_not_n841 (n841, not_n841);
	BUFX2 g_n1459 (and_pi096_pi138, n1459);
	BUFX2 g_n1558 (and_not_n1556_not_n1557, n1558);
	INVX1 g_not_pi053_4 (pi053, not_pi053_4);
	BUFX2 g_po104 (po104_driver, po104);
	BUFX2 g_n1378 (and_pi139_n1325, n1378);
	AND2X1 g_and_pi137_not_n1506 (pi137, not_n1506, and_pi137_not_n1506);
	BUFX2 g_n571 (and_n569_n570, n571);
	BUFX2 g_po127 (po127_driver, po127);
	AND2X1 g_and_not_pi024_4_not_pi042_2 (not_pi024_4, not_pi042_2, and_not_pi024_4_not_pi042_2);
	BUFX2 g_po046_driver (and_not_pi129_797922662976120010_not_n873, po046_driver);
	BUFX2 g_n604 (and_pi017_not_pi054_70, n604);
	INVX1 g_not_pi144 (pi144, not_pi144);
	BUFX2 g_n774 (and_not_pi058_0_n773, n774);
	BUFX2 g_n593 (and_not_n578_n592, n593);
	INVX1 g_not_n919 (n919, not_n919);
	BUFX2 g_po034 (po034_driver, po034);
	AND2X1 g_and_not_n1000_not_n1003 (not_n1003, not_n1000, and_not_n1000_not_n1003);
	INVX1 g_not_n979 (n979, not_n979);
	INVX1 g_not_n1232 (n1232, not_n1232);
	BUFX2 g_n1413 (and_pi138_n1246, n1413);
	INVX1 g_not_pi100 (pi100, not_pi100);
	AND2X1 g_and_pi082_not_n1027 (not_n1027, pi082, and_pi082_not_n1027);
	BUFX2 g_n831 (and_not_pi096_2_n830, n831);
	INVX1 g_not_n1197 (n1197, not_n1197);
	INVX1 g_not_n732 (n732, not_n732);
	AND2X1 g_and_n934_n1074 (n934, n1074, and_n934_n1074);
	BUFX2 g_n1229 (and_n1223_n1228, n1229);
	INVX1 g_not_n1262 (n1262, not_n1262);
	AND2X1 g_and_not_pi011_0_not_pi012_1 (not_pi012_1, not_pi011_0, and_not_pi011_0_not_pi012_1);
	INVX1 g_not_pi005_0 (pi005, not_pi005_0);
	AND2X1 g_and_pi082_not_n645 (not_n645, pi082, and_pi082_not_n645);
	BUFX2 g_po082_driver (or_pi129_n1278, po082_driver);
	AND2X1 g_and_n384_n1054 (n1054, n384, and_n384_n1054);
	AND2X1 g_and_n1251_n1281 (n1251, n1281, and_n1251_n1281);
	BUFX2 g_n1609 (and_not_pi129_1181813865805958799768684143120019644340385488367699234582870392070_not_n1608, n1609);
	BUFX2 g_n1339 (and_pi145_n1325, n1339);
	INVX1 g_not_pi003_2824752490 (pi003, not_pi003_2824752490);
	AND2X1 g_and_not_pi129_8272697060641711598380789001840137510382698418573894642080092744490_not_n1616 (not_pi129_8272697060641711598380789001840137510382698418573894642080092744490, not_n1616, and_not_pi129_8272697060641711598380789001840137510382698418573894642080092744490_not_n1616);
	INVX1 g_not_n885 (n885, not_n885);
	BUFX2 g_n971 (and_n404_n970, n971);
	BUFX2 g_po137 (po137_driver, po137);
	BUFX2 g_po056_driver (and_not_n969_n981, po056_driver);
	BUFX2 g_n1342 (and_pi082_not_n1325_3, n1342);
	INVX1 g_not_n696 (n696, not_n696);
	AND2X1 g_and_not_pi096_n714 (n714, not_pi096, and_not_pi096_n714);
	AND2X1 g_and_not_pi145_0_n1271 (n1271, not_pi145_0, and_not_pi145_0_n1271);
	AND2X1 g_and_pi010_not_pi054_5 (not_pi054_5, pi010, and_pi010_not_pi054_5);
	INVX1 g_not_n353 (n353, not_n353);
	INVX1 g_not_n719 (n719, not_n719);
	INVX1 g_not_pi085_9 (pi085, not_pi085_9);
	INVX1 g_not_pi003_273687473400809163430 (pi003, not_pi003_273687473400809163430);
	BUFX2 g_n805 (and_not_pi027_6_not_n804, n805);
	BUFX2 g_n365 (and_not_pi013_3_not_n364, n365);
	INVX1 g_not_pi002 (pi002, not_pi002);
	AND2X1 g_and_pi082_not_n391 (not_n391, pi082, and_pi082_not_n391);
	BUFX2 g_n1155 (and_n754_n1154, n1155);
	INVX1 g_not_n1144 (n1144, not_n1144);
	AND2X1 g_and_pi114_not_pi122 (not_pi122, pi114, and_pi114_not_pi122);
	INVX1 g_not_pi058 (pi058, not_pi058);
	AND2X1 g_and_not_n511_not_n519 (not_n511, not_n519, and_not_n511_not_n519);
	BUFX2 g_n1603 (and_not_n1601_not_n1602, n1603);
	BUFX2 g_po004 (po004_driver, po004);
	BUFX2 g_n659 (and_not_n657_not_n658, n659);
	BUFX2 g_n844 (and_n838_n843, n844);
	AND2X1 g_and_n408_n1088 (n408, n1088, and_n408_n1088);
	AND2X1 g_and_not_n1181_not_n1183 (not_n1183, not_n1181, and_not_n1181_not_n1183);
	AND2X1 g_and_not_n896_not_n900 (not_n896, not_n900, and_not_n896_not_n900);
	INVX1 g_not_pi011_0 (pi011, not_pi011_0);
	AND2X1 g_and_not_pi129_968890104070_not_n709 (not_n709, not_pi129_968890104070, and_not_pi129_968890104070_not_n709);
	INVX1 g_not_n530 (n530, not_n530);
	AND2X1 g_and_not_pi000_not_n306 (not_pi000, not_n306, and_not_pi000_not_n306);
	BUFX2 g_n1241 (and_not_pi122_1_n1240, n1241);
	INVX1 g_not_n1377 (n1377, not_n1377);
	AND2X1 g_and_not_pi129_185621159210175743024531636712070_not_n1096 (not_pi129_185621159210175743024531636712070, not_n1096, and_not_pi129_185621159210175743024531636712070_not_n1096);
	AND2X1 g_and_not_n1613_not_n1615 (not_n1615, not_n1613, and_not_n1613_not_n1615);
	AND2X1 g_and_not_pi129_24118650322570587750381309043265707027354805885055086420058579430_not_n1597 (not_pi129_24118650322570587750381309043265707027354805885055086420058579430, not_n1597, and_not_pi129_24118650322570587750381309043265707027354805885055086420058579430_not_n1597);
	INVX1 g_not_pi085_1 (pi085, not_pi085_1);
	INVX1 g_not_pi003_24010 (pi003, not_pi003_24010);
	INVX1 g_not_n764 (n764, not_n764);
	AND2X1 g_and_not_pi085_8_n787 (not_pi085_8, n787, and_not_pi085_8_n787);
	BUFX2 g_n649 (and_not_pi050_1_n403, n649);
	BUFX2 g_n714 (and_not_pi085_not_pi110, n714);
	AND2X1 g_and_n314_n326 (n314, n326, and_n314_n326);
	BUFX2 g_n574 (and_not_pi015_0_n573, n574);
	BUFX2 g_n504 (and_not_pi009_2_n449, n504);
	BUFX2 g_n829 (and_pi029_pi110, n829);
	INVX1 g_not_n1446 (n1446, not_n1446);
	INVX1 g_not_pi027_70 (pi027, not_pi027_70);
	BUFX2 g_n675 (and_n503_n674, n675);
	INVX1 g_not_pi120 (pi120, not_pi120);
	INVX1 g_not_n1349 (n1349, not_n1349);
	BUFX2 g_n630 (and_not_pi004_1_not_pi018_3, n630);
	INVX1 g_not_n358 (n358, not_n358);
	INVX1 g_not_pi129_1176490 (pi129, not_pi129_1176490);
	BUFX2 g_po100_driver (and_not_pi026_168070_n1375, po100_driver);
	BUFX2 g_n632 (and_n448_n631, n632);
	INVX1 g_not_n1181 (n1181, not_n1181);
	INVX1 g_not_pi007_6 (pi007, not_pi007_6);
	AND2X1 g_and_not_n793_not_n797 (not_n797, not_n793, and_not_n793_not_n797);
	BUFX2 g_po138_driver (or_pi129_pi135, po138_driver);
	AND2X1 g_and_not_pi085_0_not_n732 (not_pi085_0, not_n732, and_not_pi085_0_not_n732);
	BUFX2 g_n777 (and_pi027_pi116, n777);
	INVX1 g_not_n844 (n844, not_n844);
	BUFX2 g_n1296 (and_not_pi145_n1249, n1296);
	BUFX2 g_n1471 (and_pi034_pi136, n1471);
	INVX1 g_not_n657 (n657, not_n657);
	BUFX2 g_po117 (po117_driver, po117);
	AND2X1 g_and_not_pi026_70_pi058 (not_pi026_70, pi058, and_not_pi026_70_pi058);
	INVX1 g_not_pi009 (pi009, not_pi009);
	INVX1 g_not_n1019 (n1019, not_n1019);
	AND2X1 g_and_pi007_n357 (pi007, n357, and_pi007_n357);
	BUFX2 g_n1403 (and_pi092_not_n1386_3, n1403);
	BUFX2 g_n973 (and_pi082_not_n972, n973);
	BUFX2 g_n1217 (and_not_n1215_not_n1216, n1217);
	OR2X1 g_or_pi129_n1274 (pi129, n1274, or_pi129_n1274);
	AND2X1 g_and_pi053_not_pi085_2 (pi053, not_pi085_2, and_pi053_not_pi085_2);
	INVX1 g_not_n1386_4 (n1386, not_n1386_4);
	AND2X1 g_and_not_n368_not_n370 (not_n368, not_n370, and_not_n368_not_n370);
	BUFX2 g_po110_driver (and_not_pi129_12197604876358357001385738625629718207556152941312384010_not_n1426, po110_driver);
	BUFX2 g_n565 (and_not_n557_not_n564, n565);
	BUFX2 g_n1350 (and_pi119_pi138, n1350);
	INVX1 g_not_n1108 (n1108, not_n1108);
	AND2X1 g_and_n549_n1614 (n549, n1614, and_n549_n1614);
	INVX1 g_not_pi029_1 (pi029, not_pi029_1);
	AND2X1 g_and_not_pi026_3430_not_pi053_7 (not_pi053_7, not_pi026_3430, and_not_pi026_3430_not_pi053_7);
	BUFX2 g_po098 (po098_driver, po098);
	BUFX2 g_n551 (and_not_pi007_7_n417, n551);
	INVX1 g_not_n1070 (n1070, not_n1070);
	INVX1 g_not_pi019_0 (pi019, not_pi019_0);
	INVX1 g_not_n745 (n745, not_n745);
	INVX1 g_not_n986 (n986, not_n986);
	INVX1 g_not_n1247_2 (n1247, not_n1247_2);
	INVX1 g_not_pi110 (pi110, not_pi110);
	INVX1 g_not_n1545 (n1545, not_n1545);
	AND2X1 g_and_not_pi003_1_n470 (not_pi003_1, n470, and_not_pi003_1_n470);
	BUFX2 g_n391 (and_not_pi040_n390, n391);
	AND2X1 g_and_pi082_not_n1127 (not_n1127, pi082, and_pi082_not_n1127);
	INVX1 g_not_n1229 (n1229, not_n1229);
	AND2X1 g_and_not_pi137_not_pi138 (not_pi137, not_pi138, and_not_pi137_not_pi138);
	AND2X1 g_and_not_n1326_not_n1327 (not_n1327, not_n1326, and_not_n1326_not_n1327);
	AND2X1 g_and_pi096_pi138 (pi096, pi138, and_pi096_pi138);
	BUFX2 g_po073_driver (and_not_pi085_70_n1212, po073_driver);
	AND2X1 g_and_n408_n927 (n408, n927, and_n408_n927);
	INVX1 g_not_n1005 (n1005, not_n1005);
	BUFX2 g_n518 (and_n515_n517, n518);
	BUFX2 g_n336 (and_not_n309_not_n335, n336);
	AND2X1 g_and_not_pi144_n1249 (n1249, not_pi144, and_not_pi144_n1249);
	INVX1 g_not_n1455 (n1455, not_n1455);
	INVX1 g_not_n1102 (n1102, not_n1102);
	INVX1 g_not_n1336 (n1336, not_n1336);
	AND2X1 g_and_not_pi116_10_not_n1214 (not_pi116_10, not_n1214, and_not_pi116_10_not_n1214);
	INVX1 g_not_n1096 (n1096, not_n1096);
	INVX1 g_not_pi003_7 (pi003, not_pi003_7);
	INVX1 g_not_n625 (n625, not_n625);
	BUFX2 g_n1336 (and_not_n1334_not_n1335, n1336);
	BUFX2 g_po024_driver (and_not_pi003_4_n509, po024_driver);
	INVX1 g_not_pi017_1 (pi017, not_pi017_1);
	INVX1 g_not_n903 (n903, not_n903);
	BUFX2 g_n1455 (and_pi136_not_n1454, n1455);
	BUFX2 g_n1365 (and_pi084_not_n1325_4, n1365);
	INVX1 g_not_n1426 (n1426, not_n1426);
	BUFX2 g_n1457 (and_not_pi137_4_not_n1456, n1457);
	INVX1 g_not_pi109_4 (pi109, not_pi109_4);
	AND2X1 g_and_not_pi129_3445521474652941107197329863323672432479257983579298060008368490_n1592 (not_pi129_3445521474652941107197329863323672432479257983579298060008368490, n1592, and_not_pi129_3445521474652941107197329863323672432479257983579298060008368490_n1592);
	BUFX2 g_n1441 (and_pi141_n1386, n1441);
	BUFX2 g_n925 (and_not_pi002_2_not_pi048_2, n925);
	INVX1 g_not_n781 (n781, not_n781);
	BUFX2 g_n1200 (and_pi057_not_pi058_9, n1200);
	BUFX2 g_n1585 (and_not_n1580_not_n1584, n1585);
	INVX1 g_not_n821 (n821, not_n821);
	INVX1 g_not_n1121 (n1121, not_n1121);
	INVX1 g_not_pi003_8235430 (pi003, not_pi003_8235430);
	BUFX2 g_po062_driver (and_not_n1068_n1078, po062_driver);
	INVX1 g_not_pi016_2 (pi016, not_pi016_2);
	INVX1 g_not_pi054_9 (pi054, not_pi054_9);
	INVX1 g_not_pi003_138412872010 (pi003, not_pi003_138412872010);
	AND2X1 g_and_pi062_n1091 (n1091, pi062, and_pi062_n1091);
	INVX1 g_not_n1169 (n1169, not_n1169);
	AND2X1 g_and_not_pi043_0_n407 (not_pi043_0, n407, and_not_pi043_0_n407);
	INVX1 g_not_pi027_7 (pi027, not_pi027_7);
	INVX1 g_not_n1076 (n1076, not_n1076);
	INVX1 g_not_pi115 (pi115, not_pi115);
	AND2X1 g_and_not_n379_9_not_n1038 (not_n1038, not_n379_9, and_not_n379_9_not_n1038);
	INVX1 g_not_pi129_93874803376477543056490 (pi129, not_pi129_93874803376477543056490);
	BUFX2 g_n851 (and_pi085_n774, n851);
	AND2X1 g_and_not_pi051_1_pi109 (not_pi051_1, pi109, and_not_pi051_1_pi109);
	AND2X1 g_and_n927_n984 (n984, n927, and_n927_n984);
	BUFX2 g_po124 (po124_driver, po124);
	INVX1 g_not_n959 (n959, not_n959);
	AND2X1 g_and_n444_n445 (n444, n445, and_n444_n445);
	AND2X1 g_and_not_pi046_1_n388 (n388, not_pi046_1, and_not_pi046_1_n388);
	AND2X1 g_and_not_pi009_1_not_pi014_3 (not_pi009_1, not_pi014_3, and_not_pi009_1_not_pi014_3);
	BUFX2 g_n1075 (and_n934_n1074, n1075);
	BUFX2 g_po086_driver (or_pi129_n1298, po086_driver);
	INVX1 g_not_n829 (n829, not_n829);
	INVX1 g_not_n302 (n302, not_n302);
	INVX1 g_not_pi042_1 (pi042, not_pi042_1);
	AND2X1 g_and_not_pi137_8_not_n1519 (not_n1519, not_pi137_8, and_not_pi137_8_not_n1519);
	INVX1 g_not_n328 (n328, not_n328);
	BUFX2 g_n654 (and_pi020_not_n653, n654);
	BUFX2 g_n461 (and_not_pi028_n460, n461);
	BUFX2 g_n854 (and_not_pi026_9_not_n853, n854);
	AND2X1 g_and_not_pi002_2_not_pi048_2 (not_pi048_2, not_pi002_2, and_not_pi002_2_not_pi048_2);
	INVX1 g_not_n1285 (n1285, not_n1285);
	BUFX2 g_n1041 (and_not_pi038_2_n641, n1041);
	BUFX2 g_n1071 (and_not_n379_70_not_n1070, n1071);
	AND2X1 g_and_not_pi141_0_n1271 (n1271, not_pi141_0, and_not_pi141_0_n1271);
	AND2X1 g_and_pi082_not_n692 (pi082, not_n692, and_pi082_not_n692);
	BUFX2 g_n683 (and_not_pi129_19773267430_not_n682, n683);
	BUFX2 g_n419 (and_not_pi008_2_not_pi017_2, n419);
	BUFX2 g_n1564 (and_not_n1562_not_n1563, n1564);
	AND2X1 g_and_not_pi074_not_pi136_9 (not_pi074, not_pi136_9, and_not_pi074_not_pi136_9);
	INVX1 g_not_n1476 (n1476, not_n1476);
	AND2X1 g_and_not_n1316_not_n1317 (not_n1317, not_n1316, and_not_n1316_not_n1317);
	BUFX2 g_n1502 (and_not_n1500_not_n1501, n1502);
	BUFX2 g_po036 (po036_driver, po036);
	AND2X1 g_and_n354_n373 (n373, n354, and_n354_n373);
	AND2X1 g_and_not_pi043_3_not_n1004 (not_n1004, not_pi043_3, and_not_pi043_3_not_n1004);
	AND2X1 g_and_not_pi141_n1249 (n1249, not_pi141, and_not_pi141_n1249);
	BUFX2 g_n835 (and_not_n829_not_n834, n835);
	INVX1 g_not_pi116_7 (pi116, not_pi116_7);
	AND2X1 g_and_n441_n443 (n441, n443, and_n441_n443);
	BUFX2 g_n1191 (and_not_pi058_8_not_n1190, n1191);
	AND2X1 g_and_n583_n587 (n587, n583, and_n583_n587);
	BUFX2 g_n564 (and_n560_n563, n564);
	AND2X1 g_and_pi020_not_n653 (pi020, not_n653, and_pi020_not_n653);
	BUFX2 g_n954 (and_n388_n390, n954);
	AND2X1 g_and_n754_n1154 (n1154, n754, and_n754_n1154);
	AND2X1 g_and_not_n737_n795 (n795, not_n737, and_not_n737_n795);
	AND2X1 g_and_n1583_n1588 (n1588, n1583, and_n1583_n1588);
	BUFX2 g_n1171 (and_not_n1164_0_not_n1170, n1171);
	AND2X1 g_and_pi053_not_pi058_4 (not_pi058_4, pi053, and_pi053_not_pi058_4);
	AND2X1 g_and_not_pi142_n1249 (n1249, not_pi142, and_not_pi142_n1249);
	INVX1 g_not_n1184 (n1184, not_n1184);
	BUFX2 g_n890 (and_pi033_pi109, n890);
	BUFX2 g_n1318 (and_not_n1316_not_n1317, n1318);
	AND2X1 g_and_not_pi003_4_n509 (not_pi003_4, n509, and_not_pi003_4_n509);
	BUFX2 g_n293 (and_n291_n292, n293);
	BUFX2 g_n321 (and_not_pi014_0_not_n320, n321);
	BUFX2 g_n590 (and_pi082_not_n589, n590);
	AND2X1 g_and_pi089_pi138 (pi138, pi089, and_pi089_pi138);
	INVX1 g_not_n1397 (n1397, not_n1397);
	BUFX2 g_po084 (po084_driver, po084);
	BUFX2 g_n1017 (and_n638_n642, n1017);
	BUFX2 g_n528 (and_n416_n527, n528);
	INVX1 g_not_n1432 (n1432, not_n1432);
	BUFX2 g_n966 (and_pi082_not_n948, n966);
	INVX1 g_not_pi129_8272697060641711598380789001840137510382698418573894642080092744490 (pi129, not_pi129_8272697060641711598380789001840137510382698418573894642080092744490);
	INVX1 g_not_pi002_4 (pi002, not_pi002_4);
	BUFX2 g_n747 (and_pi025_not_pi026_1, n747);
	INVX1 g_not_pi053 (pi053, not_pi053);
	INVX1 g_not_pi129_797922662976120010 (pi129, not_pi129_797922662976120010);
	INVX1 g_not_pi146_0 (pi146, not_pi146_0);
	INVX1 g_not_pi070_0 (pi070, not_pi070_0);
	INVX1 g_not_pi138_3430 (pi138, not_pi138_3430);
	AND2X1 g_and_pi082_not_n920 (pi082, not_n920, and_pi082_not_n920);
	AND2X1 g_and_pi081_pi120 (pi120, pi081, and_pi081_pi120);
	INVX1 g_not_pi026_490 (pi026, not_pi026_490);
	BUFX2 g_n1228 (and_pi027_n1182, n1228);
	INVX1 g_not_pi136_403536070 (pi136, not_pi136_403536070);
	INVX1 g_not_n1365 (n1365, not_n1365);
	INVX1 g_not_pi007_9 (pi007, not_pi007_9);
	BUFX2 g_n1064 (and_pi082_not_n408, n1064);
	INVX1 g_not_n1452 (n1452, not_n1452);
	BUFX2 g_n459 (and_not_pi005_3_not_pi007_5, n459);
	INVX1 g_not_pi123 (pi123, not_pi123);
	BUFX2 g_n460 (and_pi025_not_pi029_0, n460);
	AND2X1 g_and_n571_n574 (n574, n571, and_n571_n574);
	BUFX2 g_n1581 (and_not_pi136_57648010_pi139, n1581);
	INVX1 g_not_n930 (n930, not_n930);
	BUFX2 g_n1080 (and_n638_n1027, n1080);
	BUFX2 g_po035 (po035_driver, po035);
	BUFX2 g_n941 (and_n736_n940, n941);
	INVX1 g_not_n1580 (n1580, not_n1580);
	BUFX2 g_n755 (and_not_pi053_0_pi058, n755);
	INVX1 g_not_n1225 (n1225, not_n1225);
	AND2X1 g_and_not_n1503_not_n1507 (not_n1503, not_n1507, and_not_n1503_not_n1507);
	BUFX2 g_n610 (and_not_pi016_2_n351, n610);
	BUFX2 g_n454 (and_n446_n453, n454);
	AND2X1 g_and_n297_n304 (n304, n297, and_n297_n304);
	AND2X1 g_and_not_pi003_9_n566 (n566, not_pi003_9, and_not_pi003_9_n566);
	INVX1 g_not_n407 (n407, not_n407);
	INVX1 g_not_n880 (n880, not_n880);
	AND2X1 g_and_pi142_n1414 (pi142, n1414, and_pi142_n1414);
	AND2X1 g_and_pi023_pi138 (pi138, pi023, and_pi023_pi138);
	AND2X1 g_and_not_pi012_3_n449 (not_pi012_3, n449, and_not_pi012_3_n449);
	BUFX2 g_n332 (and_not_pi006_0_not_pi012_0, n332);
	BUFX2 g_n352 (and_not_n350_n351, n352);
	BUFX2 g_n870 (and_pi031_not_pi109_0, n870);
	INVX1 g_not_n1114 (n1114, not_n1114);
	AND2X1 g_and_not_n691_not_n694 (not_n691, not_n694, and_not_n691_not_n694);
	INVX1 g_not_n869 (n869, not_n869);
	AND2X1 g_and_n407_n580 (n580, n407, and_n407_n580);
	BUFX2 g_po111_driver (and_not_pi129_85383234134508499009700170379408027452893070589186688070_not_n1430, po111_driver);
	BUFX2 g_n308 (and_n301_not_n302, n308);
	INVX1 g_not_n753 (n753, not_n753);
	INVX1 g_not_n1366 (n1366, not_n1366);
	AND2X1 g_and_not_n869_not_n870 (not_n870, not_n869, and_not_n869_not_n870);
	BUFX2 g_n1208 (and_n737_n1207, n1208);
	AND2X1 g_and_not_pi044_3_n379 (n379, not_pi044_3, and_not_pi044_3_n379);
	INVX1 g_not_n1414 (n1414, not_n1414);
	INVX1 g_not_pi006_2 (pi006, not_pi006_2);
	INVX1 g_not_pi003_8 (pi003, not_pi003_8);
	BUFX2 g_n381 (and_not_pi043_not_pi047, n381);
	BUFX2 g_n761 (and_pi085_not_pi116_1, n761);
	BUFX2 g_n905 (and_pi036_not_pi109_5, n905);
	BUFX2 g_po042 (po042_driver, po042);
	AND2X1 g_and_pi094_not_n1414 (pi094, not_n1414, and_pi094_not_n1414);
	AND2X1 g_and_not_n959_n962 (not_n959, n962, and_not_n959_n962);
	INVX1 g_not_pi003_0 (pi003, not_pi003_0);
	BUFX2 g_n394 (and_n386_n393, n394);
	BUFX2 g_n591 (and_pi015_n411, n591);
	BUFX2 g_n1237 (and_pi060_not_n1236, n1237);
	AND2X1 g_and_not_n379_168070_not_n1158 (not_n1158, not_n379_168070, and_not_n379_168070_not_n1158);
	BUFX2 g_n819 (and_not_pi116_4_n818, n819);
	BUFX2 g_n1517 (and_not_n1515_not_n1516, n1517);
	INVX1 g_not_pi025 (pi025, not_pi025);
	INVX1 g_not_n761 (n761, not_n761);
	INVX1 g_not_n1531 (n1531, not_n1531);
	AND2X1 g_and_not_pi137_6_not_n1491 (not_n1491, not_pi137_6, and_not_pi137_6_not_n1491);
	BUFX2 g_po108_driver (and_not_pi129_248930711762415449007872216849586085868492917169640490_not_n1409, po108_driver);
	AND2X1 g_and_not_pi038_0_not_pi040_0 (not_pi040_0, not_pi038_0, and_not_pi038_0_not_pi040_0);
	BUFX2 g_n425 (and_not_n423_n424, n425);
	AND2X1 g_and_pi138_not_n1498 (pi138, not_n1498, and_pi138_not_n1498);
	BUFX2 g_n817 (and_not_pi053_3_not_n816, n817);
	BUFX2 g_n1388 (and_pi139_n1386, n1388);
	AND2X1 g_and_not_n1458_not_n1462 (not_n1458, not_n1462, and_not_n1458_not_n1462);
	INVX1 g_not_pi085_6 (pi085, not_pi085_6);
	AND2X1 g_and_pi100_not_n716 (not_n716, pi100, and_pi100_not_n716);
	INVX1 g_not_n498 (n498, not_n498);
	BUFX2 g_n1074 (and_pi047_n641, n1074);
	BUFX2 g_n1335 (and_pi144_n1325, n1335);
	BUFX2 g_n1608 (and_n1606_n1607, n1608);
	INVX1 g_not_n1459 (n1459, not_n1459);
	OR2X1 g_or_not_pi122_2_pi129 (pi129, not_pi122_2, or_not_pi122_2_pi129);
	AND2X1 g_and_not_pi070_n577 (n577, not_pi070, and_not_pi070_n577);
	BUFX2 g_po128 (po128_driver, po128);
	INVX1 g_not_n1555 (n1555, not_n1555);
	INVX1 g_not_n469 (n469, not_n469);
	AND2X1 g_and_n1246_not_n1603 (n1246, not_n1603, and_n1246_not_n1603);
	OR2X1 g_or_n1499_n1509 (n1499, n1509, or_n1499_n1509);
	INVX1 g_not_pi041 (pi041, not_pi041);
	INVX1 g_not_pi011_2 (pi011, not_pi011_2);
	AND2X1 g_and_not_n1415_not_n1416 (not_n1416, not_n1415, and_not_n1415_not_n1416);
	AND2X1 g_and_pi079_not_n1325_0 (not_n1325_0, pi079, and_pi079_not_n1325_0);
	INVX1 g_not_pi041_0 (pi041, not_pi041_0);
	BUFX2 g_n1463 (and_not_n1458_not_n1462, n1463);
	INVX1 g_not_n1058 (n1058, not_n1058);
	AND2X1 g_and_n404_n638 (n404, n638, and_n404_n638);
	BUFX2 g_n1550 (and_pi137_not_n1549, n1550);
	BUFX2 g_n840 (and_pi058_not_n839, n840);
	BUFX2 g_n980 (and_not_pi129_225393402906922580878632490_not_n979, n980);
	INVX1 g_not_n1530 (n1530, not_n1530);
	BUFX2 g_n474 (and_pi008_not_pi017_3, n474);
	INVX1 g_not_pi028_0 (pi028, not_pi028_0);
	AND2X1 g_and_not_n379_6_not_n993 (not_n379_6, not_n993, and_not_n379_6_not_n993);
	BUFX2 g_n1604 (and_n1246_not_n1603, n1604);
	BUFX2 g_po012_driver (tie1, po012_driver);
	BUFX2 g_n1387 (and_pi088_not_n1386, n1387);
	INVX1 g_not_pi129_57908879424491981188665523012880962572678888930017262494560649211430 (pi129, not_pi129_57908879424491981188665523012880962572678888930017262494560649211430);
	AND2X1 g_and_not_pi002_0_not_pi020_0 (not_pi002_0, not_pi020_0, and_not_pi002_0_not_pi020_0);
	INVX1 g_not_n589 (n589, not_n589);
	AND2X1 g_and_pi029_not_pi116_5 (pi029, not_pi116_5, and_pi029_not_pi116_5);
	AND2X1 g_and_pi035_n1360 (n1360, pi035, and_pi035_n1360);
	AND2X1 g_and_not_n995_n997 (n997, not_n995, and_not_n995_n997);
	BUFX2 g_n887 (and_not_n882_not_n886, n887);
	INVX1 g_not_n1271_5 (n1271, not_n1271_5);
	INVX1 g_not_pi129_24010 (pi129, not_pi129_24010);
	INVX1 g_not_pi027_4 (pi027, not_pi027_4);
	AND2X1 g_and_pi082_not_n956 (not_n956, pi082, and_pi082_not_n956);
	INVX1 g_not_pi047 (pi047, not_pi047);
	INVX1 g_not_pi014 (pi014, not_pi014);
	INVX1 g_not_pi129_103677930763188441902487387275962551382129494864490 (pi129, not_pi129_103677930763188441902487387275962551382129494864490);
	BUFX2 g_n1267 (and_n1251_n1266, n1267);
	INVX1 g_not_n397 (n397, not_n397);
	AND2X1 g_and_pi137_not_n1487 (pi137, not_n1487, and_pi137_not_n1487);
	BUFX2 g_n1114 (and_pi082_not_n1113, n1114);
	BUFX2 g_n960 (and_pi040_pi082, n960);
	BUFX2 g_n959 (and_pi073_n958, n959);
	INVX1 g_not_n1260 (n1260, not_n1260);
	AND2X1 g_and_not_n1265_not_n1267 (not_n1265, not_n1267, and_not_n1265_not_n1267);
	INVX1 g_not_n1475 (n1475, not_n1475);
	INVX1 g_not_pi085 (pi085, not_pi085);
	INVX1 g_not_pi011_5 (pi011, not_pi011_5);
	INVX1 g_not_n1325_1 (n1325, not_n1325_1);
	BUFX2 g_n1338 (and_pi081_not_n1325_2, n1338);
	BUFX2 g_n855 (and_n754_n787, n855);
	AND2X1 g_and_n570_n579 (n570, n579, and_n570_n579);
	AND2X1 g_and_not_n1144_not_n1147 (not_n1147, not_n1144, and_not_n1144_not_n1147);
	INVX1 g_not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490 (pi129, not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490);
	AND2X1 g_and_n399_n568 (n399, n568, and_n399_n568);
	BUFX2 g_n516 (and_not_pi009_3_not_pi022_2, n516);
	AND2X1 g_and_not_pi129_3430_not_n565 (not_n565, not_pi129_3430, and_not_pi129_3430_not_n565);
	AND2X1 g_and_n380_n688 (n688, n380, and_n380_n688);
	AND2X1 g_and_n379_not_n1122 (n379, not_n1122, and_n379_not_n1122);
	BUFX2 g_n411 (and_not_pi082_n379, n411);
	AND2X1 g_and_not_n911_not_n912 (not_n912, not_n911, and_not_n911_not_n912);
	BUFX2 g_n1266 (and_not_pi146_n1249, n1266);
	AND2X1 g_and_not_pi042_not_pi044 (not_pi044, not_pi042, and_not_pi042_not_pi044);
	AND2X1 g_and_not_n1199_not_n1201 (not_n1201, not_n1199, and_not_n1199_not_n1201);
	AND2X1 g_and_pi013_not_pi054_8 (not_pi054_8, pi013, and_pi013_not_pi054_8);
	AND2X1 g_and_n547_n552 (n552, n547, and_n547_n552);
	INVX1 g_not_n694 (n694, not_n694);
	AND2X1 g_and_n388_n641 (n388, n641, and_n388_n641);
	INVX1 g_not_pi129_205005145156954906122290109080958673914396262484637238056070 (pi129, not_pi129_205005145156954906122290109080958673914396262484637238056070);
	INVX1 g_not_pi069 (pi069, not_pi069);
	BUFX2 g_n1133 (and_not_pi129_9095436801298611408202050198891430_not_n1132, n1133);
	INVX1 g_not_n871 (n871, not_n871);
	INVX1 g_not_pi129_70316764788835532799945507414768825152637918032230572653232010 (pi129, not_pi129_70316764788835532799945507414768825152637918032230572653232010);
	AND2X1 g_and_pi136_not_pi137_0 (not_pi137_0, pi136, and_pi136_not_pi137_0);
	BUFX2 g_n1268 (and_not_n1265_not_n1267, n1268);
	BUFX2 g_n301 (and_not_pi005_not_pi022, n301);
	INVX1 g_not_pi044_0 (pi044, not_pi044_0);
	AND2X1 g_and_not_n1334_not_n1335 (not_n1334, not_n1335, and_not_n1334_not_n1335);
	BUFX2 g_n1059 (and_pi046_pi082, n1059);
	AND2X1 g_and_pi075_n1057 (pi075, n1057, and_pi075_n1057);
	INVX1 g_not_pi138_1 (pi138, not_pi138_1);
	BUFX2 g_n1582 (and_not_pi137_70_pi138, n1582);
	BUFX2 g_n807 (and_not_n805_not_n806, n807);
	AND2X1 g_and_n1251_n1256 (n1251, n1256, and_n1251_n1256);
	INVX1 g_not_n1417 (n1417, not_n1417);
	AND2X1 g_and_n640_n644 (n640, n644, and_n640_n644);
	INVX1 g_not_n367 (n367, not_n367);
	AND2X1 g_and_not_pi061_not_pi118 (not_pi118, not_pi061, and_not_pi061_not_pi118);
	BUFX2 g_n1201 (and_n1192_n1200, n1201);
	BUFX2 g_n1530 (and_not_pi027_3430_n1529, n1530);
	BUFX2 g_n713 (and_pi085_pi116, n713);
	INVX1 g_not_n1566 (n1566, not_n1566);
	AND2X1 g_and_not_pi008_0_not_pi021_0 (not_pi021_0, not_pi008_0, and_not_pi008_0_not_pi021_0);
	INVX1 g_not_pi100_0 (pi100, not_pi100_0);
	BUFX2 g_n1092 (and_pi062_n1091, n1092);
	BUFX2 g_n772 (and_not_pi003_8235430_n771, n772);
	BUFX2 g_n1409 (and_not_n1407_not_n1408, n1409);
	INVX1 g_not_n395 (n395, not_n395);
	INVX1 g_not_pi136_57648010 (pi136, not_pi136_57648010);
	INVX1 g_not_pi047_3 (pi047, not_pi047_3);
	INVX1 g_not_n1130 (n1130, not_n1130);
	AND2X1 g_and_not_pi140_0_n1271 (n1271, not_pi140_0, and_not_pi140_0_n1271);
	AND2X1 g_and_not_pi129_19773267430_not_n682 (not_pi129_19773267430, not_n682, and_not_pi129_19773267430_not_n682);
	BUFX2 g_n550 (and_n357_n549, n550);
	AND2X1 g_and_not_pi026_490_pi037 (pi037, not_pi026_490, and_not_pi026_490_pi037);
	AND2X1 g_and_not_n1565_not_n1566 (not_n1565, not_n1566, and_not_n1565_not_n1566);
	BUFX2 g_n852 (and_n838_n851, n852);
	AND2X1 g_and_n976_n978 (n978, n976, and_n976_n978);
	INVX1 g_not_n780 (n780, not_n780);
	AND2X1 g_and_n312_n357 (n312, n357, and_n312_n357);
	AND2X1 g_and_not_n1295_not_n1297 (not_n1295, not_n1297, and_not_n1295_not_n1297);
	AND2X1 g_and_not_pi072_not_pi138_2 (not_pi138_2, not_pi072, and_not_pi072_not_pi138_2);
	BUFX2 g_po043 (po043_driver, po043);
	BUFX2 g_po087_driver (or_pi129_n1302, po087_driver);
	AND2X1 g_and_not_pi003_57648010_n785 (not_pi003_57648010, n785, and_not_pi003_57648010_n785);
	AND2X1 g_and_n927_n991 (n991, n927, and_n927_n991);
	BUFX2 g_n1220 (and_pi096_n1219, n1220);
	INVX1 g_not_pi129_1181813865805958799768684143120019644340385488367699234582870392070 (pi129, not_pi129_1181813865805958799768684143120019644340385488367699234582870392070);
	INVX1 g_not_n1064 (n1064, not_n1064);
	INVX1 g_not_pi020 (pi020, not_pi020);
	BUFX2 g_n467 (and_n447_n466, n467);
	AND2X1 g_and_not_pi018_1_not_pi021_2 (not_pi021_2, not_pi018_1, and_not_pi018_1_not_pi021_2);
	AND2X1 g_and_n294_n355 (n294, n355, and_n294_n355);
	AND2X1 g_and_not_pi003_16284135979104490_n1532 (n1532, not_pi003_16284135979104490, and_not_pi003_16284135979104490_n1532);
	AND2X1 g_and_not_pi106_9_not_n943_0 (not_pi106_9, not_n943_0, and_not_pi106_9_not_n943_0);
	INVX1 g_not_n662 (n662, not_n662);
	INVX1 g_not_pi129_225393402906922580878632490 (pi129, not_pi129_225393402906922580878632490);
	INVX1 g_not_pi129_6 (pi129, not_pi129_6);
	BUFX2 g_n769 (and_pi026_n768, n769);
	INVX1 g_not_n968 (n968, not_n968);
	BUFX2 g_n1010 (and_pi077_n1009, n1010);
	AND2X1 g_and_n381_n387 (n381, n387, and_n381_n387);
	INVX1 g_not_n379_3430 (n379, not_n379_3430);
	BUFX2 g_n1214 (and_not_n755_not_n843, n1214);
	INVX1 g_not_pi138_8235430 (pi138, not_pi138_8235430);
	BUFX2 g_po021 (po021_driver, po021);
	BUFX2 g_n1436 (and_pi098_not_n1386_5, n1436);
	BUFX2 g_n530 (and_n526_n529, n530);
	BUFX2 g_n681 (and_n675_n680, n681);
	INVX1 g_not_n879 (n879, not_n879);
	AND2X1 g_and_not_n1320_not_n1321 (not_n1320, not_n1321, and_not_n1320_not_n1321);
	AND2X1 g_and_not_n1029_not_n1032 (not_n1029, not_n1032, and_not_n1029_not_n1032);
	BUFX2 g_n782 (and_not_pi100_0_not_n781, n782);
	INVX1 g_not_n972 (n972, not_n972);
	AND2X1 g_and_not_n620_not_n624 (not_n624, not_n620, and_not_n620_not_n624);
	BUFX2 g_n988 (and_not_n983_not_n987, n988);
	INVX1 g_not_n739 (n739, not_n739);
	BUFX2 g_po034_driver (and_not_pi003_3430_n636, po034_driver);
	BUFX2 g_po006 (po006_driver, po006);
	BUFX2 g_n1514 (and_pi136_not_n1513, n1514);
	INVX1 g_not_n1391 (n1391, not_n1391);
	AND2X1 g_and_not_pi067_not_pi138_57648010 (not_pi067, not_pi138_57648010, and_not_pi067_not_pi138_57648010);
	AND2X1 g_and_not_pi047_0_not_pi048_0 (not_pi048_0, not_pi047_0, and_not_pi047_0_not_pi048_0);
	BUFX2 g_n949 (and_n389_n948, n949);
	AND2X1 g_and_not_n1150_not_n1151 (not_n1151, not_n1150, and_not_n1150_not_n1151);
	BUFX2 g_n1282 (and_n1251_n1281, n1282);
	AND2X1 g_and_pi137_not_n1567 (pi137, not_n1567, and_pi137_not_n1567);
	AND2X1 g_and_n677_n679 (n677, n679, and_n677_n679);
	INVX1 g_not_n1124 (n1124, not_n1124);
	AND2X1 g_and_not_n1178_not_n1179 (not_n1179, not_n1178, and_not_n1178_not_n1179);
	AND2X1 g_and_not_n1485_not_n1486 (not_n1486, not_n1485, and_not_n1485_not_n1486);
	BUFX2 g_n1277 (and_not_pi139_0_n1271, n1277);
	INVX1 g_not_n701 (n701, not_n701);
	AND2X1 g_and_not_pi041_2_not_n968 (not_n968, not_pi041_2, and_not_pi041_2_not_n968);
	BUFX2 g_n926 (and_n398_n925, n926);
	OR2X1 g_or_n1484_n1494 (n1494, n1484, or_n1484_n1494);
	INVX1 g_not_n1021 (n1021, not_n1021);
	INVX1 g_not_pi129_881247870897231951843937366879128181133112010 (pi129, not_pi129_881247870897231951843937366879128181133112010);
	BUFX2 g_n374 (and_n354_n373, n374);
	BUFX2 g_n555 (and_not_pi129_490_not_n554, n555);
	BUFX2 g_n317 (and_pi008_pi021, n317);
	INVX1 g_not_pi074 (pi074, not_pi074);
	INVX1 g_not_pi126 (pi126, not_pi126);
	INVX1 g_not_pi054_3 (pi054, not_pi054_3);
	BUFX2 g_n424 (and_not_pi061_not_pi118, n424);
	BUFX2 g_n602 (and_not_pi129_168070_not_n601, n602);
	AND2X1 g_and_not_pi053_0_pi058 (not_pi053_0, pi058, and_not_pi053_0_pi058);
	BUFX2 g_n765 (and_not_pi026_2_n713, n765);
	INVX1 g_not_pi022 (pi022, not_pi022);
	BUFX2 g_n876 (and_pi031_pi109, n876);
	INVX1 g_not_pi010_2 (pi010, not_pi010_2);
	BUFX2 g_po007_driver (pi101, po007_driver);
	BUFX2 g_n815 (and_n813_n814, n815);
	INVX1 g_not_n728 (n728, not_n728);
	AND2X1 g_and_n322_n516 (n516, n322, and_n322_n516);
	INVX1 g_not_n531 (n531, not_n531);
	INVX1 g_not_n716 (n716, not_n716);
	INVX1 g_not_n878 (n878, not_n878);
	INVX1 g_not_n927 (n927, not_n927);
	AND2X1 g_and_not_pi010_0_not_pi022_0 (not_pi022_0, not_pi010_0, and_not_pi010_0_not_pi022_0);
	BUFX2 g_po080_driver (or_pi129_n1268, po080_driver);
	AND2X1 g_and_not_pi129_14811132966169777414641055325137507340304213552070_not_n1389 (not_n1389, not_pi129_14811132966169777414641055325137507340304213552070, and_not_pi129_14811132966169777414641055325137507340304213552070_not_n1389);
	INVX1 g_not_n604 (n604, not_n604);
	OR2X1 g_or_pi129_n1310 (n1310, pi129, or_pi129_n1310);
	XNOR2X1 g_tie1 (pi048, pi048, tie1);
	INVX1 g_not_pi011_3 (pi011, not_pi011_3);
	AND2X1 g_and_not_pi139_0_n1271 (n1271, not_pi139_0, and_not_pi139_0_n1271);
	BUFX2 g_n722 (and_not_pi051_not_pi052, n722);
	INVX1 g_not_n1378 (n1378, not_n1378);
	AND2X1 g_and_pi016_not_pi054_10 (pi016, not_pi054_10, and_pi016_not_pi054_10);
	BUFX2 g_n1067 (and_not_n1064_not_n1066, n1067);
	INVX1 g_not_n1436 (n1436, not_n1436);
	BUFX2 g_n1234 (and_not_pi129_7490483309651862334944941026945644936490_not_n1233, n1234);
	AND2X1 g_and_not_pi129_85383234134508499009700170379408027452893070589186688070_not_n1430 (not_pi129_85383234134508499009700170379408027452893070589186688070, not_n1430, and_not_pi129_85383234134508499009700170379408027452893070589186688070_not_n1430);
	INVX1 g_not_n1030 (n1030, not_n1030);
	AND2X1 g_and_n384_n586 (n586, n384, and_n384_n586);
	BUFX2 g_n666 (and_n299_n665, n666);
	INVX1 g_not_n1556 (n1556, not_n1556);
	BUFX2 g_n1221 (and_not_n1218_not_n1220, n1221);
	INVX1 g_not_n1450 (n1450, not_n1450);
	AND2X1 g_and_not_n1034_n1046 (not_n1034, n1046, and_not_n1034_n1046);
	AND2X1 g_and_not_n1005_n1015 (n1015, not_n1005, and_not_n1005_n1015);
	INVX1 g_not_pi116_8 (pi116, not_pi116_8);
	AND2X1 g_and_not_pi001_not_n352 (not_n352, not_pi001, and_not_pi001_not_n352);
	INVX1 g_not_n799 (n799, not_n799);
	BUFX2 g_n1150 (and_pi097_n1149, n1150);
	INVX1 g_not_n983 (n983, not_n983);
	BUFX2 g_n1511 (and_pi092_pi138, n1511);
	INVX1 g_not_n363 (n363, not_n363);
	AND2X1 g_and_n385_n698 (n385, n698, and_n385_n698);
	BUFX2 g_n670 (and_not_pi129_2824752490_not_n669, n670);
	INVX1 g_not_n1090 (n1090, not_n1090);
	AND2X1 g_and_pi082_not_n1055 (pi082, not_n1055, and_pi082_not_n1055);
	BUFX2 g_n502 (and_n499_n501, n502);
	AND2X1 g_and_pi065_not_n1247_2 (pi065, not_n1247_2, and_pi065_not_n1247_2);
	BUFX2 g_n658 (and_pi020_n411, n658);
	BUFX2 g_n1395 (and_pi090_not_n1386_1, n1395);
	INVX1 g_not_pi085_490 (pi085, not_pi085_490);
	INVX1 g_not_pi106_2 (pi106, not_pi106_2);
	BUFX2 g_n729 (and_not_n727_not_n728, n729);
	INVX1 g_not_po129 (po129_driver, not_po129);
	AND2X1 g_and_not_pi129_26517308458596534717790233816010_not_n1076 (not_pi129_26517308458596534717790233816010, not_n1076, and_not_pi129_26517308458596534717790233816010_not_n1076);
	INVX1 g_not_n394 (n394, not_n394);
	AND2X1 g_and_pi044_pi082 (pi044, pi082, and_pi044_pi082);
	BUFX2 g_n1442 (and_not_n1440_not_n1441, n1442);
	BUFX2 g_n1244 (and_pi136_n1243, n1244);
	BUFX2 g_n865 (and_pi088_pi106, n865);
	OR2X1 g_or_pi129_pi134 (pi129, pi134, or_pi129_pi134);
	INVX1 g_not_n1280 (n1280, not_n1280);
	AND2X1 g_and_pi092_not_n1386_3 (not_n1386_3, pi092, and_pi092_not_n1386_3);
	BUFX2 g_po005_driver (pi105, po005_driver);
	INVX1 g_not_pi007_5 (pi007, not_pi007_5);
	INVX1 g_not_n482 (n482, not_n482);
	AND2X1 g_and_n450_n610 (n610, n450, and_n450_n610);
	BUFX2 g_po080 (po080_driver, po080);
	AND2X1 g_and_pi082_not_n985 (not_n985, pi082, and_pi082_not_n985);
	BUFX2 g_po026_driver (and_not_pi003_6_n532, po026_driver);
	BUFX2 g_n357 (and_not_pi005_1_n332, n357);
	INVX1 g_not_pi007 (pi007, not_pi007);
	INVX1 g_not_n410 (n410, not_n410);
	AND2X1 g_and_n927_n929 (n929, n927, and_n927_n929);
	AND2X1 g_and_not_n940_not_n1136 (not_n1136, not_n940, and_not_n940_not_n1136);
	BUFX2 g_po101 (po101_driver, po101);
	BUFX2 g_po083_driver (or_pi129_n1283, po083_driver);
	BUFX2 g_n1021 (and_not_pi044_3_n379, n1021);
	BUFX2 g_n736 (and_not_pi039_0_not_pi052_0, n736);
	INVX1 g_not_n576 (n576, not_n576);
	BUFX2 g_n794 (and_pi026_not_pi027_5, n794);
	AND2X1 g_and_pi074_n932 (n932, pi074, and_pi074_n932);
	AND2X1 g_and_not_n1349_not_n1353 (not_n1353, not_n1349, and_not_n1349_not_n1353);
	AND2X1 g_and_not_pi010_not_n324 (not_n324, not_pi010, and_not_pi010_not_n324);
	INVX1 g_not_n472 (n472, not_n472);
	AND2X1 g_and_not_pi028_0_n548 (n548, not_pi028_0, and_not_pi028_0_n548);
	INVX1 g_not_n1173 (n1173, not_n1173);
	BUFX2 g_n1298 (and_not_n1295_not_n1297, n1298);
	BUFX2 g_n1081 (and_pi082_not_n1080, n1081);
	INVX1 g_not_pi110_5 (pi110, not_pi110_5);
	INVX1 g_not_n1405 (n1405, not_n1405);
	BUFX2 g_n693 (and_pi082_not_n692, n693);
	BUFX2 g_n1072 (and_pi064_n1071, n1072);
	BUFX2 g_n382 (and_n380_n381, n382);
	AND2X1 g_and_not_pi085_6_not_n849 (not_pi085_6, not_n849, and_not_pi085_6_not_n849);
	BUFX2 g_n994 (and_not_n379_6_not_n993, n994);
	BUFX2 g_n620 (and_pi018_not_pi054_490, n620);
	AND2X1 g_and_pi054_not_pi059_0 (not_pi059_0, pi054, and_pi054_not_pi059_0);
	INVX1 g_not_n922 (n922, not_n922);
	BUFX2 g_po113_driver (and_not_pi129_4183778472590916451475308348590993345191760458870147715430_not_n1438, po113_driver);
	AND2X1 g_and_not_n379_5_not_n973 (not_n973, not_n379_5, and_not_n379_5_not_n973);
	AND2X1 g_and_n918_n1043 (n1043, n918, and_n918_n1043);
	INVX1 g_not_pi003_6782230728490 (pi003, not_pi003_6782230728490);
	INVX1 g_not_n1308 (n1308, not_n1308);
	BUFX2 g_n969 (and_not_pi041_2_not_n968, n969);
	AND2X1 g_and_not_n969_n981 (n981, not_n969, and_not_n969_n981);
	BUFX2 g_n294 (and_not_pi017_not_pi021, n294);
	AND2X1 g_and_n1087_n1120 (n1120, n1087, and_n1087_n1120);
	INVX1 g_not_pi058_0 (pi058, not_pi058_0);
	BUFX2 g_n1596 (and_pi054_not_n1595, n1596);
	BUFX2 g_po062 (po062_driver, po062);
	INVX1 g_not_pi116_3 (pi116, not_pi116_3);
	INVX1 g_not_n884 (n884, not_n884);
	INVX1 g_not_n379_10 (n379, not_n379_10);
	AND2X1 g_and_pi063_not_n1247_0 (not_n1247_0, pi063, and_pi063_not_n1247_0);
	BUFX2 g_n1487 (and_not_n1485_not_n1486, n1487);
	BUFX2 g_n315 (and_pi007_not_n311, n315);
	BUFX2 g_po122 (po122_driver, po122);
	INVX1 g_not_n794_0 (n794, not_n794_0);
	BUFX2 g_n430 (and_pi010_not_pi022_1, n430);
	INVX1 g_not_n1471 (n1471, not_n1471);
	AND2X1 g_and_n419_n473 (n473, n419, and_n419_n473);
	BUFX2 g_n801 (and_not_pi110_2_n800, n801);
	INVX1 g_not_n1596 (n1596, not_n1596);
	INVX1 g_not_n311 (n311, not_n311);
	INVX1 g_not_n656 (n656, not_n656);
	INVX1 g_not_n908 (n908, not_n908);
	AND2X1 g_and_not_n425_not_n427 (not_n427, not_n425, and_not_n425_not_n427);
	INVX1 g_not_pi069_0 (pi069, not_pi069_0);
	OR2X1 g_or_pi123_pi129 (pi129, pi123, or_pi123_pi129);
	AND2X1 g_and_n536_n537 (n537, n536, and_n536_n537);
	AND2X1 g_and_pi030_not_pi109 (pi030, not_pi109, and_pi030_not_pi109);
	AND2X1 g_and_pi082_not_n949 (not_n949, pi082, and_pi082_not_n949);
	INVX1 g_not_pi138_70 (pi138, not_pi138_70);
	BUFX2 g_n579 (and_not_pi048_1_n381, n579);
	BUFX2 g_n1314 (and_not_n1312_not_n1313, n1314);
	BUFX2 g_n1358 (and_not_n1356_not_n1357, n1358);
	BUFX2 g_n542 (and_not_pi129_70_not_n541, n542);
	INVX1 g_not_n742 (n742, not_n742);
	INVX1 g_not_pi129_113988951853731430 (pi129, not_pi129_113988951853731430);
	AND2X1 g_and_pi026_pi116 (pi116, pi026, and_pi026_pi116);
	BUFX2 g_po123 (po123_driver, po123);
	INVX1 g_not_pi095 (pi095, not_pi095);
	AND2X1 g_and_pi082_not_n394 (not_n394, pi082, and_pi082_not_n394);
	BUFX2 g_n784 (and_not_n782_not_n783, n784);
	INVX1 g_not_n1470 (n1470, not_n1470);
	AND2X1 g_and_not_pi027_6_not_n804 (not_n804, not_pi027_6, and_not_pi027_6_not_n804);
	AND2X1 g_and_not_pi136_2824752490_pi140 (not_pi136_2824752490, pi140, and_not_pi136_2824752490_pi140);
	INVX1 g_not_pi043 (pi043, not_pi043);
	AND2X1 g_and_not_pi044_0_n401 (n401, not_pi044_0, and_not_pi044_0_n401);
	INVX1 g_not_n861 (n861, not_n861);
	BUFX2 g_po058_driver (and_not_n1005_n1015, po058_driver);
	INVX1 g_not_pi004_2 (pi004, not_pi004_2);
	AND2X1 g_and_not_pi129_168070_not_n601 (not_pi129_168070, not_n601, and_not_pi129_168070_not_n601);
	INVX1 g_not_pi110_6 (pi110, not_pi110_6);
	AND2X1 g_and_n383_n384 (n383, n384, and_n383_n384);
	INVX1 g_not_n795 (n795, not_n795);
	AND2X1 g_and_n404_n406 (n406, n404, and_n404_n406);
	BUFX2 g_n1086 (and_not_pi002_4_not_pi047_4, n1086);
	BUFX2 g_n1126 (and_n404_n638, n1126);
	BUFX2 g_n1182 (and_not_pi085_8_n787, n1182);
	AND2X1 g_and_not_pi129_8_not_n508 (not_n508, not_pi129_8, and_not_pi129_8_not_n508);
	BUFX2 g_n541 (and_not_n534_not_n540, n541);
	INVX1 g_not_n1344 (n1344, not_n1344);
	AND2X1 g_and_pi002_n645 (pi002, n645, and_pi002_n645);
	AND2X1 g_and_n1246_not_n1421 (n1246, not_n1421, and_n1246_not_n1421);
	AND2X1 g_and_not_pi085_3430_not_n725_0 (not_n725_0, not_pi085_3430, and_not_pi085_3430_not_n725_0);
	BUFX2 g_po003_driver (pi103, po003_driver);
	AND2X1 g_and_pi033_pi109 (pi033, pi109, and_pi033_pi109);
	BUFX2 g_n1505 (and_pi032_pi136, n1505);
	BUFX2 g_n323 (and_n314_n322, n323);
	BUFX2 g_n492 (and_n448_n491, n492);
	INVX1 g_not_pi026_70 (pi026, not_pi026_70);
	AND2X1 g_and_pi008_not_pi054_3 (not_pi054_3, pi008, and_pi008_not_pi054_3);
	AND2X1 g_and_not_pi040_2_not_n952 (not_n952, not_pi040_2, and_not_pi040_2_not_n952);
	INVX1 g_not_n391 (n391, not_n391);
	INVX1 g_not_n914 (n914, not_n914);
	BUFX2 g_n1602 (and_not_pi115_0_not_n1421_2, n1602);
	AND2X1 g_and_not_pi022_3_n449 (not_pi022_3, n449, and_not_pi022_3_n449);
	BUFX2 g_n685 (and_not_pi023_pi055, n685);
	BUFX2 g_n810 (and_pi028_not_pi116_3, n810);
	BUFX2 g_n449 (and_not_pi004_0_not_pi019_0, n449);
	INVX1 g_not_pi109 (pi109, not_pi109);
	BUFX2 g_n409 (and_n402_n408, n409);
	BUFX2 g_n1084 (and_not_n1081_not_n1083, n1084);
	INVX1 g_not_n333 (n333, not_n333);
	AND2X1 g_and_not_pi010_2_pi022 (not_pi010_2, pi022, and_not_pi010_2_pi022);
	AND2X1 g_and_n927_n1126 (n927, n1126, and_n927_n1126);
	BUFX2 g_n1568 (and_pi137_not_n1567, n1568);
	INVX1 g_not_n1127 (n1127, not_n1127);
	BUFX2 g_po019_driver (and_not_pi003_n438, po019_driver);
	INVX1 g_not_n845 (n845, not_n845);
	BUFX2 g_n1205 (and_n814_n1169, n1205);
	INVX1 g_not_n653 (n653, not_n653);
	AND2X1 g_and_pi035_not_pi109_4 (not_pi109_4, pi035, and_pi035_not_pi109_4);
	BUFX2 g_n742 (and_not_n740_not_n741, n742);
	BUFX2 g_n299 (and_not_pi004_not_pi016, n299);
	AND2X1 g_and_n814_n1169 (n814, n1169, and_n814_n1169);
	AND2X1 g_and_not_pi050_2_n391 (n391, not_pi050_2, and_not_pi050_2_n391);
	BUFX2 g_n951 (and_n379_not_n950, n951);
	BUFX2 g_n469 (and_not_n458_not_n468, n469);
	INVX1 g_not_pi045_2 (pi045, not_pi045_2);
	BUFX2 g_po102_driver (and_not_pi129_2115876138024253916377293617876786762900601936010_not_n1383, po102_driver);
	AND2X1 g_and_not_pi003_1176490_n759 (not_pi003_1176490, n759, and_not_pi003_1176490_n759);
	INVX1 g_not_n840 (n840, not_n840);
	INVX1 g_not_pi109_0 (pi109, not_pi109_0);
	BUFX2 g_n499 (and_n291_n344, n499);
	AND2X1 g_and_n638_n1110 (n638, n1110, and_n638_n1110);
	AND2X1 g_and_not_pi129_1176490_not_n617 (not_n617, not_pi129_1176490, and_not_pi129_1176490_not_n617);
	AND2X1 g_and_n934_n1094 (n934, n1094, and_n934_n1094);
	INVX1 g_not_n634 (n634, not_n634);
	INVX1 g_not_pi043_0 (pi043, not_pi043_0);
	BUFX2 g_n1589 (and_n1583_n1588, n1589);
	INVX1 g_not_pi027_3 (pi027, not_pi027_3);
	INVX1 g_not_n1271_0 (n1271, not_n1271_0);
	BUFX2 g_n1044 (and_n918_n1043, n1044);
	INVX1 g_not_pi003_2 (pi003, not_pi003_2);
	OR2X1 g_or_pi129_n1322 (pi129, n1322, or_pi129_n1322);
	AND2X1 g_and_not_n472_not_n482 (not_n472, not_n482, and_not_n472_not_n482);
	AND2X1 g_and_n490_n492 (n492, n490, and_n490_n492);
	AND2X1 g_and_not_n350_n351 (not_n350, n351, and_not_n350_n351);
	AND2X1 g_and_n381_n406 (n406, n381, and_n381_n406);
	BUFX2 g_n405 (and_not_pi046_0_not_pi050_0, n405);
	BUFX2 g_n1371 (and_pi096_n1370, n1371);
	INVX1 g_not_pi041_1 (pi041, not_pi041_1);
	BUFX2 g_n417 (and_n344_n416, n417);
	AND2X1 g_and_pi033_pi136 (pi033, pi136, and_pi033_pi136);
	BUFX2 g_n746 (and_not_pi053_not_n745, n746);
	BUFX2 g_n566 (and_not_pi129_3430_not_n565, n566);
	BUFX2 g_n1222 (and_not_pi085_490_not_n1221, n1222);
	BUFX2 g_n1451 (and_not_pi136_4_not_n1450, n1451);
	AND2X1 g_and_pi145_n1414 (n1414, pi145, and_pi145_n1414);
	INVX1 g_not_pi039_0 (pi039, not_pi039_0);
	BUFX2 g_n1238 (and_pi123_n1236, n1238);
	INVX1 g_not_n1271_4 (n1271, not_n1271_4);
	INVX1 g_not_n792 (n792, not_n792);
	INVX1 g_not_n1478 (n1478, not_n1478);
	INVX1 g_not_n1265 (n1265, not_n1265);
	BUFX2 g_n1467 (and_pi095_n1324, n1467);
	BUFX2 g_n331 (and_not_pi017_0_n330, n331);
	BUFX2 g_n768 (and_not_pi085_4_not_n738_0, n768);
	BUFX2 g_n1301 (and_not_pi140_0_n1271, n1301);
	BUFX2 g_n1353 (and_not_pi136_1_not_n1352, n1353);
	INVX1 g_not_n737 (n737, not_n737);
	BUFX2 g_n617 (and_not_n604_not_n616, n617);
	BUFX2 g_n1096 (and_n1093_n1095, n1096);
	INVX1 g_not_pi054_0 (pi054, not_pi054_0);
	BUFX2 g_n773 (and_not_pi027_2_not_pi053_1, n773);
	BUFX2 g_n776 (and_pi095_not_pi096_1, n776);
	INVX1 g_not_pi008_2 (pi008, not_pi008_2);
	BUFX2 g_po037_driver (and_not_pi003_168070_n683, po037_driver);
	BUFX2 g_n745 (and_not_n735_not_n744, n745);
	AND2X1 g_and_pi006_not_pi012_4 (pi006, not_pi012_4, and_pi006_not_pi012_4);
	BUFX2 g_po057 (po057_driver, po057);
	AND2X1 g_and_n1246_not_n1585 (n1246, not_n1585, and_n1246_not_n1585);
	AND2X1 g_and_pi137_not_n1362 (pi137, not_n1362, and_pi137_not_n1362);
	BUFX2 g_n1065 (and_pi082_not_n927, n1065);
	AND2X1 g_and_not_pi143_0_n1249 (n1249, not_pi143_0, and_not_pi143_0_n1249);
	AND2X1 g_and_not_pi014_2_pi054 (not_pi014_2, pi054, and_not_pi014_2_pi054);
	INVX1 g_not_n915 (n915, not_n915);
	BUFX2 g_n1042 (and_pi045_n1041, n1042);
	BUFX2 g_po103_driver (and_not_pi129_14811132966169777414641055325137507340304213552070_not_n1389, po103_driver);
	BUFX2 g_n837 (and_pi097_pi116, n837);
	BUFX2 g_n1121 (and_n1087_n1120, n1121);
	BUFX2 g_po029 (po029_driver, po029);
	INVX1 g_not_n1615 (n1615, not_n1615);
	INVX1 g_not_n1191 (n1191, not_n1191);
	BUFX2 g_n892 (and_not_n890_not_n891, n892);
	BUFX2 g_n1561 (and_not_pi137_10_not_n1560, n1561);
	BUFX2 g_po094_driver (and_not_pi129_2569235775210588780886114772242356213216070_not_n1332, po094_driver);
	BUFX2 g_po055 (po055_driver, po055);
	AND2X1 g_and_not_pi129_11044276742439206463052992010_not_n1013 (not_pi129_11044276742439206463052992010, not_n1013, and_not_pi129_11044276742439206463052992010_not_n1013);
	BUFX2 g_n1223 (and_pi059_not_pi116_70, n1223);
	AND2X1 g_and_not_pi071_n647 (n647, not_pi071, and_not_pi071_n647);
	INVX1 g_not_n1233 (n1233, not_n1233);
	INVX1 g_not_n858 (n858, not_n858);
	BUFX2 g_n396 (and_not_n379_not_n395, n396);
	BUFX2 g_n453 (and_n447_n452, n453);
	BUFX2 g_n1033 (and_not_n1029_not_n1032, n1033);
	AND2X1 g_and_not_n836_not_n840 (not_n840, not_n836, and_not_n836_not_n840);
	AND2X1 g_and_not_pi013_1_pi014 (pi014, not_pi013_1, and_not_pi013_1_pi014);
	BUFX2 g_n588 (and_n583_n587, n588);
	BUFX2 g_n1559 (and_not_pi136_1176490_not_n1558, n1559);
	BUFX2 g_po050 (po050_driver, po050);
	INVX1 g_not_n726_0 (n726, not_n726_0);
	INVX1 g_not_n853 (n853, not_n853);
	INVX1 g_not_pi109_1 (pi109, not_pi109_1);
	AND2X1 g_and_n379_not_n1065 (n379, not_n1065, and_n379_not_n1065);
	BUFX2 g_n1165 (and_pi026_not_pi058_6, n1165);
	AND2X1 g_and_not_pi122_1_n1240 (n1240, not_pi122_1, and_not_pi122_1_n1240);
	INVX1 g_not_pi113_0 (pi113, not_pi113_0);
	BUFX2 g_n1109 (and_not_pi002_5_n383, n1109);
	INVX1 g_not_pi110_7 (pi110, not_pi110_7);
	BUFX2 g_n1190 (and_not_n1187_not_n1189, n1190);
	BUFX2 g_n383 (and_not_pi015_not_pi020, n383);
	AND2X1 g_and_n1192_n1196 (n1192, n1196, and_n1192_n1196);
	OR2X1 g_or_n1355_n1363 (n1355, n1363, or_n1355_n1363);
	BUFX2 g_n1513 (and_not_n1511_not_n1512, n1513);
	AND2X1 g_and_pi093_not_n1386_4 (pi093, not_n1386_4, and_pi093_not_n1386_4);
	BUFX2 g_n940 (and_not_pi051_1_pi109, n940);
	AND2X1 g_and_not_pi011_3_n449 (not_pi011_3, n449, and_not_pi011_3_n449);
	AND2X1 g_and_not_n1215_not_n1216 (not_n1215, not_n1216, and_not_n1215_not_n1216);
	BUFX2 g_n1575 (and_not_pi097_1_n755, n1575);
	BUFX2 g_n1325 (and_n1251_n1324, n1325);
	AND2X1 g_and_not_n1395_not_n1396 (not_n1395, not_n1396, and_not_n1395_not_n1396);
	INVX1 g_not_pi129_1577753820348458066150427430 (pi129, not_pi129_1577753820348458066150427430);
	INVX1 g_not_pi017_2 (pi017, not_pi017_2);
	AND2X1 g_and_pi145_n1325 (n1325, pi145, and_pi145_n1325);
	BUFX2 g_n597 (and_not_pi005_5_n596, n597);
	BUFX2 g_n720 (and_not_n717_not_n719, n720);
	INVX1 g_not_pi122_2 (pi122, not_pi122_2);
	INVX1 g_not_n508 (n508, not_n508);
	INVX1 g_not_pi045_3 (pi045, not_pi045_3);
	BUFX2 g_n1327 (and_pi142_n1325, n1327);
	BUFX2 g_n1360 (and_pi136_not_pi138_4, n1360);
	INVX1 g_not_pi138_57648010 (pi138, not_pi138_57648010);
	INVX1 g_not_n1441 (n1441, not_n1441);
	AND2X1 g_and_n728_n737 (n737, n728, and_n728_n737);
	AND2X1 g_and_not_n1555_not_n1559 (not_n1559, not_n1555, and_not_n1555_not_n1559);
	BUFX2 g_n1554 (and_not_n1552_not_n1553, n1554);
	BUFX2 g_n490 (and_n488_n489, n490);
	AND2X1 g_and_pi097_pi138 (pi138, pi097, and_pi097_pi138);
	BUFX2 g_n327 (and_n314_n326, n327);
	BUFX2 g_n1381 (and_pi087_not_n1325_6, n1381);
	AND2X1 g_and_not_n721_not_n733 (not_n721, not_n733, and_not_n721_not_n733);
	BUFX2 g_n738 (and_pi116_n737, n738);
	INVX1 g_not_n1525 (n1525, not_n1525);
	BUFX2 g_n1005 (and_not_pi043_3_not_n1004, n1005);
	BUFX2 g_n822 (and_not_n817_not_n821, n822);
	BUFX2 g_n953 (and_not_pi040_2_not_n952, n953);
	INVX1 g_not_pi129_168070 (pi129, not_pi129_168070);
	BUFX2 g_n1090 (and_pi082_not_n1089, n1090);
	AND2X1 g_and_not_pi129_12197604876358357001385738625629718207556152941312384010_not_n1426 (not_pi129_12197604876358357001385738625629718207556152941312384010, not_n1426, and_not_pi129_12197604876358357001385738625629718207556152941312384010_not_n1426);
	AND2X1 g_and_n344_n374 (n344, n374, and_n344_n374);
	AND2X1 g_and_n448_n491 (n448, n491, and_n448_n491);
	INVX1 g_not_pi025_1 (pi025, not_pi025_1);
	BUFX2 g_n1230 (and_not_n1227_not_n1229, n1230);
	INVX1 g_not_n338 (n338, not_n338);
	AND2X1 g_and_not_pi129_29286449308136415160327158440136953416342323212091034008010_not_n1442 (not_pi129_29286449308136415160327158440136953416342323212091034008010, not_n1442, and_not_pi129_29286449308136415160327158440136953416342323212091034008010_not_n1442);
	BUFX2 g_n1461 (and_not_n1459_not_n1460, n1461);
	BUFX2 g_n1488 (and_pi137_not_n1487, n1488);
	AND2X1 g_and_pi081_not_pi138_1176490 (pi081, not_pi138_1176490, and_pi081_not_pi138_1176490);
	BUFX2 g_po059_driver (and_not_n1023_n1024, po059_driver);
	INVX1 g_not_pi008_1 (pi008, not_pi008_1);
	BUFX2 g_po133_driver (and_not_pi129_8272697060641711598380789001840137510382698418573894642080092744490_not_n1616, po133_driver);
	INVX1 g_not_pi003_1176490 (pi003, not_pi003_1176490);
	AND2X1 g_and_not_pi047_3_not_n1067 (not_n1067, not_pi047_3, and_not_pi047_3_not_n1067);
	INVX1 g_not_pi018_1 (pi018, not_pi018_1);
	INVX1 g_not_n891 (n891, not_n891);
	AND2X1 g_and_n404_n970 (n404, n970, and_n404_n970);
	BUFX2 g_n942 (and_not_pi106_7_not_n941, n942);
	BUFX2 g_n992 (and_n927_n991, n992);
	BUFX2 g_n1320 (and_pi077_not_n1271_6, n1320);
	AND2X1 g_and_not_n1601_not_n1602 (not_n1602, not_n1601, and_not_n1601_not_n1602);
	AND2X1 g_and_n355_n488 (n355, n488, and_n355_n488);
	INVX1 g_not_pi122 (pi122, not_pi122);
	BUFX2 g_n624 (and_n487_n623, n624);
	AND2X1 g_and_n573_n689 (n573, n689, and_n573_n689);
	AND2X1 g_and_not_n924_n938 (n938, not_n924, and_not_n924_n938);
	AND2X1 g_and_not_pi018_not_pi019 (not_pi019, not_pi018, and_not_pi018_not_pi019);
	INVX1 g_not_n798 (n798, not_n798);
	AND2X1 g_and_not_pi085_9_not_n1188 (not_pi085_9, not_n1188, and_not_pi085_9_not_n1188);
	BUFX2 g_n1243 (and_not_pi137_not_pi138, n1243);
	OR2X1 g_or_pi129_n1306 (pi129, n1306, or_pi129_n1306);
	INVX1 g_not_n757 (n757, not_n757);
	BUFX2 g_po069 (po069_driver, po069);
	AND2X1 g_and_not_pi126_pi132 (pi132, not_pi126, and_not_pi126_pi132);
	BUFX2 g_po045 (po045_driver, po045);
	INVX1 g_not_pi022_4 (pi022, not_pi022_4);
	BUFX2 g_n456 (and_not_pi129_4_not_n455, n456);
	AND2X1 g_and_n344_n416 (n344, n416, and_n344_n416);
	AND2X1 g_and_pi037_not_pi109_6 (pi037, not_pi109_6, and_pi037_not_pi109_6);
	BUFX2 g_n586 (and_n408_n585, n586);
	INVX1 g_not_pi028 (pi028, not_pi028);
	AND2X1 g_and_pi086_not_n1325_5 (not_n1325_5, pi086, and_pi086_not_n1325_5);
	AND2X1 g_and_pi054_n1610 (n1610, pi054, and_pi054_n1610);
	BUFX2 g_po059 (po059_driver, po059);
	BUFX2 g_po119_driver (or_n1499_n1509, po119_driver);
	INVX1 g_not_n1404 (n1404, not_n1404);
	BUFX2 g_po141_driver (and_pi133_n1631, po141_driver);
	AND2X1 g_and_pi036_pi109 (pi036, pi109, and_pi036_pi109);
	AND2X1 g_and_pi060_pi109 (pi060, pi109, and_pi060_pi109);
	INVX1 g_not_n573 (n573, not_n573);
	BUFX2 g_po116 (po116_driver, po116);
	BUFX2 g_n1068 (and_not_pi047_3_not_n1067, n1068);
	AND2X1 g_and_not_pi045_not_pi048 (not_pi045, not_pi048, and_not_pi045_not_pi048);
	INVX1 g_not_n1300 (n1300, not_n1300);
	AND2X1 g_and_pi048_n1041 (pi048, n1041, and_pi048_n1041);
	INVX1 g_not_pi009_4 (pi009, not_pi009_4);
	AND2X1 g_and_not_pi075_not_pi138_490 (not_pi075, not_pi138_490, and_not_pi075_not_pi138_490);
	BUFX2 g_n553 (and_n547_n552, n553);
	AND2X1 g_and_not_n1119_not_n1123 (not_n1123, not_n1119, and_not_n1119_not_n1123);
	INVX1 g_not_pi005 (pi005, not_pi005);
	BUFX2 g_n1460 (and_pi082_not_pi138_7, n1460);
	AND2X1 g_and_not_n779_not_n780 (not_n780, not_n779, and_not_n779_not_n780);
	BUFX2 g_n1493 (and_not_n1488_not_n1492, n1493);
	AND2X1 g_and_not_pi003_n438 (n438, not_pi003, and_not_pi003_n438);
	BUFX2 g_n503 (and_n419_n473, n503);
	AND2X1 g_and_n379_not_n1031 (not_n1031, n379, and_n379_not_n1031);
	BUFX2 g_n432 (and_n369_n431, n432);
	BUFX2 g_n1039 (and_not_n379_9_not_n1038, n1039);
	AND2X1 g_and_not_pi097_1_n755 (n755, not_pi097_1, and_not_pi097_1_n755);
	AND2X1 g_and_n382_n385 (n385, n382, and_n382_n385);
	BUFX2 g_n1166 (and_pi116_n1165, n1166);
	INVX1 g_not_pi129_725745515342319093317411710931737859674906464051430 (pi129, not_pi129_725745515342319093317411710931737859674906464051430);
	BUFX2 g_po054 (po054_driver, po054);
	BUFX2 g_n509 (and_not_pi129_8_not_n508, n509);
	BUFX2 g_n809 (and_not_pi085_5_not_n808, n809);
	BUFX2 g_n1592 (and_n1246_not_n1591, n1592);
	INVX1 g_not_n1342 (n1342, not_n1342);
	INVX1 g_not_n1358 (n1358, not_n1358);
	BUFX2 g_n806 (and_n777_n790, n806);
	BUFX2 g_n733 (and_not_pi085_0_not_n732, n733);
	INVX1 g_not_pi136_3430 (pi136, not_pi136_3430);
	AND2X1 g_and_n1093_n1095 (n1093, n1095, and_n1093_n1095);
	AND2X1 g_and_not_pi007_0_pi013 (pi013, not_pi007_0, and_not_pi007_0_pi013);
	BUFX2 g_n646 (and_pi082_not_n645, n646);
	BUFX2 g_po038 (po038_driver, po038);
	BUFX2 g_n1037 (and_n408_n1036, n1037);
	BUFX2 g_n1093 (and_n381_n406, n1093);
	AND2X1 g_and_n918_n919 (n919, n918, and_n918_n919);
	INVX1 g_not_n721 (n721, not_n721);
	BUFX2 g_n1631 (and_not_pi126_pi132, n1631);
	AND2X1 g_and_not_n735_not_n744 (not_n744, not_n735, and_not_n735_not_n744);
	BUFX2 g_n389 (and_n387_n388, n389);
	INVX1 g_not_pi116_10 (pi116, not_pi116_10);
	BUFX2 g_n1285 (and_pi069_not_n1247_4, n1285);
	BUFX2 g_po089 (po089_driver, po089);
	AND2X1 g_and_n381_n405 (n405, n381, and_n381_n405);
	BUFX2 g_n1088 (and_n1086_n1087, n1088);
	INVX1 g_not_n1267 (n1267, not_n1267);
	INVX1 g_not_n1052 (n1052, not_n1052);
	BUFX2 g_n752 (and_not_n746_not_n751, n752);
	BUFX2 g_n1422 (and_n1246_not_n1421, n1422);
	AND2X1 g_and_not_pi136_0_pi137 (pi137, not_pi136_0, and_not_pi136_0_pi137);
	AND2X1 g_and_not_pi021_3_pi054 (not_pi021_3, pi054, and_not_pi021_3_pi054);
	AND2X1 g_and_not_n1514_not_n1518 (not_n1518, not_n1514, and_not_n1514_not_n1518);
	AND2X1 g_and_n448_n504 (n448, n504, and_n448_n504);
	INVX1 g_not_n812 (n812, not_n812);
	BUFX2 g_n489 (and_not_pi011_2_pi021, n489);
	BUFX2 g_n1273 (and_not_pi143_n1271, n1273);
	INVX1 g_not_n1629 (n1629, not_n1629);
	INVX1 g_not_n1317 (n1317, not_n1317);
	AND2X1 g_and_not_n523_not_n530 (not_n530, not_n523, and_not_n523_not_n530);
	INVX1 g_not_n805 (n805, not_n805);
	BUFX2 g_n369 (and_n345_n357, n369);
	AND2X1 g_and_pi082_not_n1080 (not_n1080, pi082, and_pi082_not_n1080);
	BUFX2 g_n1179 (and_n787_n1175, n1179);
	BUFX2 g_n787 (and_not_pi053_2_not_pi058_1, n787);
	BUFX2 g_n823 (and_not_pi058_2_not_n822, n823);
	INVX1 g_not_pi137_3 (pi137, not_pi137_3);
	AND2X1 g_and_not_n1544_not_n1548 (not_n1548, not_n1544, and_not_n1544_not_n1548);
	AND2X1 g_and_not_pi085_70_n1212 (n1212, not_pi085_70, and_not_pi085_70_n1212);
	AND2X1 g_and_not_pi058_10_n1206 (not_pi058_10, n1206, and_not_pi058_10_n1206);
	AND2X1 g_and_not_pi024_2_not_n695 (not_n695, not_pi024_2, and_not_pi024_2_not_n695);
	BUFX2 g_n790 (and_not_pi026_4_not_n723_0, n790);
	BUFX2 g_n575 (and_n571_n574, n575);
	INVX1 g_not_n1217 (n1217, not_n1217);
	AND2X1 g_and_n359_n361 (n361, n359, and_n359_n361);
	AND2X1 g_and_not_n1428_not_n1429 (not_n1429, not_n1428, and_not_n1428_not_n1429);
	INVX1 g_not_pi046_1 (pi046, not_pi046_1);
	INVX1 g_not_n777 (n777, not_n777);
	BUFX2 g_po054_driver (and_not_pi129_4599865365447399609768010_not_n945, po054_driver);
	INVX1 g_not_pi051_0 (pi051, not_pi051_0);
	INVX1 g_not_pi021_1 (pi021, not_pi021_1);
	AND2X1 g_and_not_pi024_0_not_pi045_0 (not_pi045_0, not_pi024_0, and_not_pi024_0_not_pi045_0);
	BUFX2 g_n576 (and_pi082_not_n575, n576);
	AND2X1 g_and_n356_n372 (n356, n372, and_n356_n372);
	BUFX2 g_n1386 (and_n1251_n1385, n1386);
	INVX1 g_not_pi003 (pi003, not_pi003);
	AND2X1 g_and_not_pi129_490_not_n554 (not_pi129_490, not_n554, and_not_pi129_490_not_n554);
	BUFX2 g_n614 (and_n612_n613, n614);
	BUFX2 g_n1408 (and_pi146_n1386, n1408);
	AND2X1 g_and_n748_n756 (n756, n748, and_n748_n756);
	BUFX2 g_n465 (and_not_pi006_2_n450, n465);
	BUFX2 g_n326 (and_pi010_n291, n326);
	AND2X1 g_and_not_pi097_n724 (n724, not_pi097, and_not_pi097_n724);
	INVX1 g_not_n315 (n315, not_n315);
	BUFX2 g_n781 (and_not_n779_not_n780, n781);
	BUFX2 g_n878 (and_not_n876_not_n877, n878);
	AND2X1 g_and_not_pi129_77309937197074445241370944070_not_n983_0 (not_n983_0, not_pi129_77309937197074445241370944070, and_not_pi129_77309937197074445241370944070_not_n983_0);
	BUFX2 g_n633 (and_n629_n632, n633);
	AND2X1 g_and_n649_n651 (n651, n649, and_n649_n651);
	BUFX2 g_n648 (and_not_pi071_n647, n648);
	BUFX2 g_n1202 (and_not_n1199_not_n1201, n1202);
	INVX1 g_not_n725_0 (n725, not_n725_0);
	INVX1 g_not_n1424 (n1424, not_n1424);
	AND2X1 g_and_not_pi014_1_n347 (not_pi014_1, n347, and_not_pi014_1_n347);
	AND2X1 g_and_not_pi025_1_not_pi028_1 (not_pi028_1, not_pi025_1, and_not_pi025_1_not_pi028_1);
	AND2X1 g_and_pi098_pi106 (pi098, pi106, and_pi098_pi106);
	BUFX2 g_n452 (and_n448_n451, n452);
	AND2X1 g_and_not_pi129_1070069044235980333563563003849377848070_not_n1209 (not_n1209, not_pi129_1070069044235980333563563003849377848070, and_not_pi129_1070069044235980333563563003849377848070_not_n1209);
	INVX1 g_not_n1421_2 (n1421, not_n1421_2);
	AND2X1 g_and_n787_n847 (n787, n847, and_n787_n847);
	AND2X1 g_and_pi145_n1386 (n1386, pi145, and_pi145_n1386);
	AND2X1 g_and_n448_n545 (n545, n448, and_n448_n545);
	INVX1 g_not_n1321 (n1321, not_n1321);
	INVX1 g_not_pi100_2 (pi100, not_pi100_2);
	AND2X1 g_and_not_pi003_490_n626 (not_pi003_490, n626, and_not_pi003_490_n626);
	BUFX2 g_n704 (and_not_pi043_2_n387, n704);
	BUFX2 g_po076 (po076_driver, po076);
	BUFX2 g_n1370 (and_not_pi110_5_n1369, n1370);
	INVX1 g_not_pi129_248930711762415449007872216849586085868492917169640490 (pi129, not_pi129_248930711762415449007872216849586085868492917169640490);
	BUFX2 g_n402 (and_n400_n401, n402);
	INVX1 g_not_n1515 (n1515, not_n1515);
	OR2X1 g_or_n1469_n1479 (n1479, n1469, or_n1469_n1479);
	AND2X1 g_and_n369_n431 (n369, n431, and_n369_n431);
	OR2X1 g_or_pi129_n1283 (n1283, pi129, or_pi129_n1283);
	BUFX2 g_n912 (and_pi037_not_pi109_6, n912);
	BUFX2 g_po053_driver (and_not_n924_n938, po053_driver);
	INVX1 g_not_pi014_3 (pi014, not_pi014_3);
	BUFX2 g_n672 (and_pi022_not_pi054_168070, n672);
	INVX1 g_not_pi027_0 (pi027, not_pi027_0);
	BUFX2 g_n1106 (and_n990_n1105, n1106);
	INVX1 g_not_n379_24010 (n379, not_n379_24010);
	BUFX2 g_n1152 (and_not_n1150_not_n1151, n1152);
	BUFX2 g_n1189 (and_not_pi085_9_not_n1188, n1189);
	BUFX2 g_n1385 (and_pi136_pi137, n1385);
	INVX1 g_not_n1522 (n1522, not_n1522);
	AND2X1 g_and_not_pi129_1435036016098684342856030763566710717400773837392460666392490_not_n1531 (not_n1531, not_pi129_1435036016098684342856030763566710717400773837392460666392490, and_not_pi129_1435036016098684342856030763566710717400773837392460666392490_not_n1531);
	AND2X1 g_and_not_pi129_57908879424491981188665523012880962572678888930017262494560649211430_not_n724 (not_n724, not_pi129_57908879424491981188665523012880962572678888930017262494560649211430, and_not_pi129_57908879424491981188665523012880962572678888930017262494560649211430_not_n724);
	AND2X1 g_and_not_pi003_10_n602 (not_pi003_10, n602, and_not_pi003_10_n602);
	AND2X1 g_and_not_pi085_5_not_n808 (not_pi085_5, not_n808, and_not_pi085_5_not_n808);
	AND2X1 g_and_not_pi044_1_pi082 (pi082, not_pi044_1, and_not_pi044_1_pi082);
	AND2X1 g_and_not_n1104_n1116 (not_n1104, n1116, and_not_n1104_n1116);
	BUFX2 g_n370 (and_pi009_n369, n370);
	BUFX2 g_n1586 (and_n1246_not_n1585, n1586);
	BUFX2 g_n1257 (and_n1251_n1256, n1257);
	INVX1 g_not_pi137_8 (pi137, not_pi137_8);
	BUFX2 g_n1496 (and_pi099_n1249, n1496);
	INVX1 g_not_pi054_8 (pi054, not_pi054_8);
	INVX1 g_not_pi136_2824752490 (pi136, not_pi136_2824752490);
	AND2X1 g_and_n1223_n1224 (n1223, n1224, and_n1223_n1224);
	BUFX2 g_po068 (po068_driver, po068);
	INVX1 g_not_pi058_6 (pi058, not_pi058_6);
	INVX1 g_not_n1466 (n1466, not_n1466);
	INVX1 g_not_pi045_0 (pi045, not_pi045_0);
	INVX1 g_not_n947 (n947, not_n947);
	INVX1 g_not_n1000 (n1000, not_n1000);
	AND2X1 g_and_not_n1556_not_n1557 (not_n1556, not_n1557, and_not_n1556_not_n1557);
	AND2X1 g_and_pi074_not_n1271_3 (not_n1271_3, pi074, and_pi074_not_n1271_3);
	INVX1 g_not_n826 (n826, not_n826);
	AND2X1 g_and_n515_n517 (n515, n517, and_n515_n517);
	BUFX2 g_n324 (and_not_n321_not_n323, n324);
	BUFX2 g_n407 (and_n404_n406, n407);
	BUFX2 g_n443 (and_pi028_n442, n443);
	AND2X1 g_and_not_n1276_not_n1277 (not_n1276, not_n1277, and_not_n1276_not_n1277);
	INVX1 g_not_pi066 (pi066, not_pi066);
	INVX1 g_not_n1188 (n1188, not_n1188);
	AND2X1 g_and_n638_n928 (n638, n928, and_n638_n928);
	BUFX2 g_po056 (po056_driver, po056);
	INVX1 g_not_n923 (n923, not_n923);
	INVX1 g_not_pi010_1 (pi010, not_pi010_1);
	INVX1 g_not_n1107 (n1107, not_n1107);
	BUFX2 g_n1425 (and_pi143_n1414, n1425);
	AND2X1 g_and_n369_n528 (n528, n369, and_n369_n528);
	AND2X1 g_and_n473_n474 (n473, n474, and_n473_n474);
	AND2X1 g_and_not_n1424_not_n1425 (not_n1424, not_n1425, and_not_n1424_not_n1425);
	BUFX2 g_n605 (and_not_pi007_8_n346, n605);
	BUFX2 g_n1098 (and_not_n1092_n1097, n1098);
	AND2X1 g_and_not_pi007_6_n449 (not_pi007_6, n449, and_not_pi007_6_n449);
	AND2X1 g_and_not_pi002_1_not_pi045_3 (not_pi045_3, not_pi002_1, and_not_pi002_1_not_pi045_3);
	BUFX2 g_n609 (and_n445_n608, n609);
	BUFX2 g_n1521 (and_pi080_not_pi138_3430, n1521);
	AND2X1 g_and_not_pi145_n1249 (n1249, not_pi145, and_not_pi145_n1249);
	BUFX2 g_n418 (and_n347_n417, n418);
	BUFX2 g_n780 (and_not_pi027_3_n713, n780);
	INVX1 g_not_pi141_0 (pi141, not_pi141_0);
	AND2X1 g_and_pi096_n1370 (pi096, n1370, and_pi096_n1370);
	BUFX2 g_n1103 (and_not_n379_3430_not_n1102, n1103);
	INVX1 g_not_n703 (n703, not_n703);
	AND2X1 g_and_not_pi136_8235430_not_n1564 (not_pi136_8235430, not_n1564, and_not_pi136_8235430_not_n1564);
	INVX1 g_not_n758 (n758, not_n758);
	BUFX2 g_n694 (and_n379_not_n693, n694);
	BUFX2 g_n1444 (and_pi100_not_n1423_2, n1444);
	INVX1 g_not_pi146 (pi146, not_pi146);
	AND2X1 g_and_not_n696_n711 (not_n696, n711, and_not_n696_n711);
	BUFX2 g_n1031 (and_pi082_not_n1030, n1031);
	BUFX2 g_n598 (and_n345_n597, n598);
	BUFX2 g_po129_driver (or_pi123_pi129, po129_driver);
	BUFX2 g_po006_driver (pi107, po006_driver);
	BUFX2 g_n519 (and_n514_n518, n519);
	BUFX2 g_n1260 (and_pi064_not_n1247_1, n1260);
	AND2X1 g_and_n402_n408 (n408, n402, and_n402_n408);
	INVX1 g_not_pi039 (pi039, not_pi039);
	AND2X1 g_and_not_n1081_not_n1083 (not_n1081, not_n1083, and_not_n1081_not_n1083);
	INVX1 g_not_n1559 (n1559, not_n1559);
	AND2X1 g_and_not_pi106_1_not_n878 (not_pi106_1, not_n878, and_not_pi106_1_not_n878);
	BUFX2 g_n726 (and_not_pi110_0_not_n725, n726);
	INVX1 g_not_n1423 (n1423, not_n1423);
	INVX1 g_not_pi049_0 (pi049, not_pi049_0);
	BUFX2 g_n1169 (and_pi058_not_pi116_7, n1169);
	BUFX2 g_n628 (and_pi019_not_pi054_3430, n628);
	BUFX2 g_n447 (and_not_pi059_n356, n447);
	INVX1 g_not_pi085_0 (pi085, not_pi085_0);
	INVX1 g_not_n1040 (n1040, not_n1040);
	BUFX2 g_n1454 (and_not_n1452_not_n1453, n1454);
	BUFX2 g_n1468 (and_not_n1466_not_n1467, n1468);
	AND2X1 g_and_not_pi068_pi136 (pi136, not_pi068, and_not_pi068_pi136);
	INVX1 g_not_n1564 (n1564, not_n1564);
	BUFX2 g_n339 (and_not_pi129_not_n338, n339);
	BUFX2 g_n967 (and_n379_not_n966, n967);
	AND2X1 g_and_pi082_not_n573 (pi082, not_n573, and_pi082_not_n573);
	INVX1 g_not_n1485 (n1485, not_n1485);
	INVX1 g_not_n1247_6 (n1247, not_n1247_6);
	AND2X1 g_and_not_pi096_2_n830 (not_pi096_2, n830, and_not_pi096_2_n830);
	BUFX2 g_po005 (po005_driver, po005);
	AND2X1 g_and_n448_n535 (n535, n448, and_n448_n535);
	INVX1 g_not_pi002_2 (pi002, not_pi002_2);
	AND2X1 g_and_n538_n539 (n539, n538, and_n538_n539);
	AND2X1 g_and_not_n578_n592 (not_n578, n592, and_not_n578_n592);
	INVX1 g_not_pi007_2 (pi007, not_pi007_2);
	AND2X1 g_and_n1054_n1059 (n1054, n1059, and_n1054_n1059);
	BUFX2 g_po109_driver (and_not_pi129_1742514982336908143055105517947102601079450420187483430_not_n1417, po109_driver);
	AND2X1 g_and_pi125_pi138 (pi125, pi138, and_pi125_pi138);
	AND2X1 g_and_pi116_n737 (n737, pi116, and_pi116_n737);
	INVX1 g_not_n336 (n336, not_n336);
	AND2X1 g_and_not_n837_not_n838 (not_n838, not_n837, and_not_n837_not_n838);
	INVX1 g_not_n941 (n941, not_n941);
	INVX1 g_not_pi009_6 (pi009, not_pi009_6);
	BUFX2 g_n1304 (and_pi073_not_n1271_2, n1304);
	INVX1 g_not_pi010_0 (pi010, not_pi010_0);
	INVX1 g_not_n943_0 (n943, not_n943_0);
	BUFX2 g_n1215 (and_not_pi116_10_not_n1214, n1215);
	AND2X1 g_and_not_n486_not_n494 (not_n486, not_n494, and_not_n486_not_n494);
	INVX1 g_not_pi100_1 (pi100, not_pi100_1);
	AND2X1 g_and_pi032_pi109 (pi032, pi109, and_pi032_pi109);
	INVX1 g_not_n591 (n591, not_n591);
	INVX1 g_not_n1423_0 (n1423, not_n1423_0);
	AND2X1 g_and_n380_n1111 (n380, n1111, and_n380_n1111);
	AND2X1 g_and_n1581_n1583 (n1581, n1583, and_n1581_n1583);
	INVX1 g_not_pi129_125892552985318850263419623839875454447587430 (pi129, not_pi129_125892552985318850263419623839875454447587430);
	BUFX2 g_n669 (and_not_n662_not_n668, n669);
	INVX1 g_not_n320 (n320, not_n320);
	BUFX2 g_n663 (and_n355_n488, n663);
	BUFX2 g_po051_driver (and_not_pi129_13410686196639649008070_not_n908, po051_driver);
	BUFX2 g_n1046 (and_not_n1040_n1045, n1046);
	BUFX2 g_po127_driver (and_not_pi129_3445521474652941107197329863323672432479257983579298060008368490_n1592, po127_driver);
	INVX1 g_not_pi006_1 (pi006, not_pi006_1);
	INVX1 g_not_pi110_0 (pi110, not_pi110_0);
	BUFX2 g_n1020 (and_pi067_not_n379_8, n1020);
	AND2X1 g_and_not_pi003_797922662976120010_n1577 (n1577, not_pi003_797922662976120010, and_not_pi003_797922662976120010_n1577);
	INVX1 g_not_pi040_2 (pi040, not_pi040_2);
	INVX1 g_not_n993 (n993, not_n993);
	INVX1 g_not_n1123 (n1123, not_n1123);
	INVX1 g_not_n685 (n685, not_n685);
	AND2X1 g_and_pi005_not_n332 (not_n332, pi005, and_pi005_not_n332);
	INVX1 g_not_pi047_4 (pi047, not_pi047_4);
	AND2X1 g_and_not_n379_not_n395 (not_n395, not_n379, and_not_n379_not_n395);
	BUFX2 g_n1506 (and_not_n1504_not_n1505, n1506);
	INVX1 g_not_pi022_2 (pi022, not_pi022_2);
	INVX1 g_not_pi129_6168735096280623662907561568153897267931784070 (pi129, not_pi129_6168735096280623662907561568153897267931784070);
	BUFX2 g_n642 (and_n388_n641, n642);
	AND2X1 g_and_n380_n381 (n380, n381, and_n380_n381);
	INVX1 g_not_pi129_367033682172941254412302110320336601888010 (pi129, not_pi129_367033682172941254412302110320336601888010);
	INVX1 g_not_n752 (n752, not_n752);
	BUFX2 g_n1501 (and_not_pi073_not_pi136_10, n1501);
	INVX1 g_not_n796 (n796, not_n796);
	INVX1 g_not_pi026_168070 (pi026, not_pi026_168070);
	BUFX2 g_n494 (and_n487_n493, n494);
	BUFX2 g_n1464 (and_pi137_not_n1463, n1464);
	INVX1 g_not_n808 (n808, not_n808);
	AND2X1 g_and_pi085_n718 (n718, pi085, and_pi085_n718);
	AND2X1 g_and_not_n854_not_n857 (not_n857, not_n854, and_not_n854_not_n857);
	INVX1 g_not_pi138_8 (pi138, not_pi138_8);
	INVX1 g_not_n1023 (n1023, not_n1023);
	INVX1 g_not_n985 (n985, not_n985);
	AND2X1 g_and_not_n868_not_n872 (not_n872, not_n868, and_not_n868_not_n872);
	INVX1 g_not_n1430 (n1430, not_n1430);
	BUFX2 g_po082 (po082_driver, po082);
	INVX1 g_not_n723 (n723, not_n723);
	BUFX2 g_n1236 (and_not_pi117_not_pi122_0, n1236);
	INVX1 g_not_n1290 (n1290, not_n1290);
	AND2X1 g_and_not_pi136_3_n1411 (not_pi136_3, n1411, and_not_pi136_3_n1411);
	BUFX2 g_po001_driver (pi083, po001_driver);
	AND2X1 g_and_not_pi007_2_not_pi013_2 (not_pi007_2, not_pi013_2, and_not_pi007_2_not_pi013_2);
	INVX1 g_not_pi003_3 (pi003, not_pi003_3);
	AND2X1 g_and_pi082_not_n992 (pi082, not_n992, and_pi082_not_n992);
	BUFX2 g_n1328 (and_not_n1326_not_n1327, n1328);
	AND2X1 g_and_pi096_n1219 (pi096, n1219, and_pi096_n1219);
	AND2X1 g_and_pi143_n1386 (n1386, pi143, and_pi143_n1386);
	BUFX2 g_n1573 (and_not_pi003_113988951853731430_n1572, n1573);
	INVX1 g_not_pi042_0 (pi042, not_pi042_0);
	INVX1 g_not_n1354 (n1354, not_n1354);
	BUFX2 g_n757 (and_n748_n756, n757);
	AND2X1 g_and_not_pi085_7_not_n1177 (not_n1177, not_pi085_7, and_not_pi085_7_not_n1177);
	BUFX2 g_n585 (and_not_pi015_1_not_n584, n585);
	AND2X1 g_and_not_n1260_not_n1262 (not_n1262, not_n1260, and_not_n1260_not_n1262);
	BUFX2 g_n889 (and_pi091_pi106, n889);
	AND2X1 g_and_not_n1488_not_n1492 (not_n1492, not_n1488, and_not_n1488_not_n1492);
	INVX1 g_not_pi003_39098210485829880490 (pi003, not_pi003_39098210485829880490);
	INVX1 g_not_n1542 (n1542, not_n1542);
	BUFX2 g_po027_driver (and_not_pi003_7_n542, po027_driver);
	AND2X1 g_and_not_n1140_n1141 (n1141, not_n1140, and_not_n1140_n1141);
	OR2X1 g_or_pi129_pi135 (pi135, pi129, or_pi129_pi135);
	BUFX2 g_po135 (po135_driver, po135);
	INVX1 g_not_pi110_2 (pi110, not_pi110_2);
	INVX1 g_not_n740 (n740, not_n740);
	BUFX2 g_n922 (and_n379_not_n921, n922);
	INVX1 g_not_n1216 (n1216, not_n1216);
	AND2X1 g_and_not_pi129_797922662976120010_not_n873 (not_pi129_797922662976120010, not_n873, and_not_pi129_797922662976120010_not_n873);
	BUFX2 g_n495 (and_not_n486_not_n494, n495);
	AND2X1 g_and_not_pi129_2326305139872070_not_n826 (not_n826, not_pi129_2326305139872070, and_not_pi129_2326305139872070_not_n826);
	BUFX2 g_n1177 (and_not_n1174_not_n1176, n1177);
	AND2X1 g_and_pi142_n1325 (n1325, pi142, and_pi142_n1325);
	AND2X1 g_and_not_pi006_2_n450 (not_pi006_2, n450, and_not_pi006_2_n450);
	INVX1 g_not_pi009_0 (pi009, not_pi009_0);
	AND2X1 g_and_n345_n346 (n346, n345, and_n345_n346);
	AND2X1 g_and_n813_n814 (n814, n813, and_n813_n814);
	AND2X1 g_and_pi077_n1009 (pi077, n1009, and_pi077_n1009);
	BUFX2 g_n1024 (and_not_pi129_77309937197074445241370944070_not_n983_0, n1024);
	BUFX2 g_n814 (and_not_pi026_7_not_pi027_7, n814);
	BUFX2 g_n1062 (and_not_n1058_n1061, n1062);
	INVX1 g_not_pi085_70 (pi085, not_pi085_70);
	INVX1 g_not_pi067 (pi067, not_pi067);
	BUFX2 g_n320 (and_not_n313_not_n319, n320);
	BUFX2 g_n334 (and_not_n310_not_n333, n334);
	AND2X1 g_and_pi038_n641 (n641, pi038, and_pi038_n641);
	BUFX2 g_n989 (and_not_pi042_1_not_n988, n989);
	BUFX2 g_po058 (po058_driver, po058);
	BUFX2 g_n380 (and_not_pi045_not_pi048, n380);
	BUFX2 g_n607 (and_not_pi012_5_n606, n607);
	AND2X1 g_and_n560_n563 (n563, n560, and_n560_n563);
	INVX1 g_not_n660 (n660, not_n660);
	BUFX2 g_n996 (and_pi042_n934, n996);
	AND2X1 g_and_pi138_not_n1483 (pi138, not_n1483, and_pi138_not_n1483);
	BUFX2 g_n481 (and_n445_n480, n481);
	BUFX2 g_n1614 (and_pi054_not_pi059_0, n1614);
	INVX1 g_not_pi027_10 (pi027, not_pi027_10);
	AND2X1 g_and_not_pi041_not_pi046 (not_pi041, not_pi046, and_not_pi041_not_pi046);
	INVX1 g_not_n1248 (n1248, not_n1248);
	BUFX2 g_n846 (and_not_pi027_9_not_n845, n846);
	BUFX2 g_po040_driver (and_not_pi003_1176490_n759, po040_driver);
	AND2X1 g_and_not_n1381_not_n1382 (not_n1382, not_n1381, and_not_n1381_not_n1382);
	AND2X1 g_and_pi093_pi138 (pi093, pi138, and_pi093_pi138);
	BUFX2 g_n441 (and_not_pi007_4_n332, n441);
	AND2X1 g_and_n688_n927 (n688, n927, and_n688_n927);
	INVX1 g_not_n1425 (n1425, not_n1425);
	AND2X1 g_and_not_pi009_3_not_pi022_2 (not_pi022_2, not_pi009_3, and_not_pi009_3_not_pi022_2);
	AND2X1 g_and_not_pi003_3_n496 (not_pi003_3, n496, and_not_pi003_3_n496);
	BUFX2 g_n696 (and_not_pi024_2_not_n695, n696);
	AND2X1 g_and_not_n713_not_n715 (not_n713, not_n715, and_not_n713_not_n715);
	BUFX2 g_n298 (and_not_pi018_not_pi019, n298);
	AND2X1 g_and_n723_n727 (n727, n723, and_n723_n727);
	INVX1 g_not_pi144_0 (pi144, not_pi144_0);
	AND2X1 g_and_not_pi004_0_not_pi019_0 (not_pi019_0, not_pi004_0, and_not_pi004_0_not_pi019_0);
	INVX1 g_not_n1359 (n1359, not_n1359);
	INVX1 g_not_pi058_4 (pi058, not_pi058_4);
	BUFX2 g_po090_driver (or_pi129_n1314, po090_driver);
	BUFX2 g_n526 (and_n503_n525, n526);
	BUFX2 g_n292 (and_not_pi006_not_pi007, n292);
	BUFX2 g_n545 (and_not_pi013_5_n450, n545);
	OR2X1 g_or_pi003_not_n377 (not_n377, pi003, or_pi003_not_n377);
	AND2X1 g_and_not_pi042_1_not_n988 (not_pi042_1, not_n988, and_not_pi042_1_not_n988);
	AND2X1 g_and_not_pi138_8_not_n1478 (not_pi138_8, not_n1478, and_not_pi138_8_not_n1478);
	BUFX2 g_n987 (and_n379_not_n986, n987);
	BUFX2 g_po072 (po072_driver, po072);
	AND2X1 g_and_not_pi137_7_not_n1502 (not_n1502, not_pi137_7, and_not_pi137_7_not_n1502);
	BUFX2 g_n375 (and_n344_n374, n375);
	BUFX2 g_n367 (and_not_n365_not_n366, n367);
	BUFX2 g_n1176 (and_not_pi058_7_n1175, n1176);
	BUFX2 g_n1052 (and_not_n1048_not_n1051, n1052);
	INVX1 g_not_n301 (n301, not_n301);
	INVX1 g_not_n454 (n454, not_n454);
	BUFX2 g_n679 (and_n479_n678, n679);
	AND2X1 g_and_not_n1280_not_n1282 (not_n1280, not_n1282, and_not_n1280_not_n1282);
	AND2X1 g_and_not_pi110_0_not_n725 (not_n725, not_pi110_0, and_not_pi110_0_not_n725);
	AND2X1 g_and_not_pi106_3_not_n892 (not_pi106_3, not_n892, and_not_pi106_3_not_n892);
	BUFX2 g_n877 (and_pi032_not_pi109_1, n877);
	INVX1 g_not_n843 (n843, not_n843);
	AND2X1 g_and_pi066_not_n1271 (pi066, not_n1271, and_pi066_not_n1271);
	BUFX2 g_n1181 (and_not_pi027_10_not_n1180, n1181);
	BUFX2 g_n483 (and_not_n472_not_n482, n483);
	INVX1 g_not_n723_0 (n723, not_n723_0);
	AND2X1 g_and_pi027_n768 (n768, pi027, and_pi027_n768);
	BUFX2 g_n923 (and_not_n917_not_n922, n923);
	INVX1 g_not_pi097_0 (pi097, not_pi097_0);
	BUFX2 g_n1619 (and_not_pi110_7_not_pi120, n1619);
	BUFX2 g_n1518 (and_not_pi136_490_not_n1517, n1518);
	BUFX2 g_n1193 (and_not_pi116_9_n1192, n1193);
	BUFX2 g_n638 (and_n381_n387, n638);
	INVX1 g_not_n1350 (n1350, not_n1350);
	INVX1 g_not_pi138_24010 (pi138, not_pi138_24010);
	BUFX2 g_n1343 (and_pi146_n1325, n1343);
	INVX1 g_not_pi007_10 (pi007, not_pi007_10);
	AND2X1 g_and_not_pi027_4_n737 (not_pi027_4, n737, and_not_pi027_4_n737);
	AND2X1 g_and_not_pi129_597682638941559493067901192655856192170251494124306816490_not_n1434 (not_pi129_597682638941559493067901192655856192170251494124306816490, not_n1434, and_not_pi129_597682638941559493067901192655856192170251494124306816490_not_n1434);
	INVX1 g_not_n428 (n428, not_n428);
	INVX1 g_not_pi027_9 (pi027, not_pi027_9);
	INVX1 g_not_n862 (n862, not_n862);
	INVX1 g_not_pi045_4 (pi045, not_pi045_4);
	AND2X1 g_and_not_pi129_1577753820348458066150427430_not_n996 (not_pi129_1577753820348458066150427430, not_n996, and_not_pi129_1577753820348458066150427430_not_n996);
	BUFX2 g_n1432 (and_pi097_not_n1423_1, n1432);
	BUFX2 g_n413 (and_pi002_not_n412, n413);
	BUFX2 g_n950 (and_pi082_not_n949, n950);
	BUFX2 g_n997 (and_not_pi129_1577753820348458066150427430_not_n996, n997);
	BUFX2 g_po039_driver (and_not_n696_n711, po039_driver);
	AND2X1 g_and_not_pi015_not_pi020 (not_pi015, not_pi020, and_not_pi015_not_pi020);
	INVX1 g_not_pi106_1 (pi106, not_pi106_1);
	INVX1 g_not_n1001 (n1001, not_n1001);
	BUFX2 g_n1565 (and_not_pi136_8235430_not_n1564, n1565);
	BUFX2 g_n883 (and_pi032_pi109, n883);
	INVX1 g_not_n1044 (n1044, not_n1044);
	BUFX2 g_po139 (po139_driver, po139);
	BUFX2 g_n1354 (and_not_n1349_not_n1353, n1354);
	AND2X1 g_and_not_pi066_not_pi136_7 (not_pi066, not_pi136_7, and_not_pi066_not_pi136_7);
	BUFX2 g_n908 (and_not_n903_not_n907, n908);
	AND2X1 g_and_n1251_n1266 (n1251, n1266, and_n1251_n1266);
	INVX1 g_not_n1158 (n1158, not_n1158);
	AND2X1 g_and_pi140_n1386 (n1386, pi140, and_pi140_n1386);
	AND2X1 g_and_pi066_n1129 (pi066, n1129, and_pi066_n1129);
	BUFX2 g_po093_driver (and_not_pi129_367033682172941254412302110320336601888010_not_n1328, po093_driver);
	INVX1 g_not_n833 (n833, not_n833);
	AND2X1 g_and_pi144_n1325 (n1325, pi144, and_pi144_n1325);
	AND2X1 g_and_not_pi003_5_n521 (n521, not_pi003_5, and_not_pi003_5_n521);
	AND2X1 g_and_n300_n342 (n342, n300, and_n300_n342);
	BUFX2 g_po086 (po086_driver, po086);
	INVX1 g_not_n857 (n857, not_n857);
	BUFX2 g_po044 (po044_driver, po044);
	INVX1 g_not_n1032 (n1032, not_n1032);
	AND2X1 g_and_pi082_not_n404 (pi082, not_n404, and_pi082_not_n404);
	INVX1 g_not_pi136_1 (pi136, not_pi136_1);
	INVX1 g_not_pi137_9 (pi137, not_pi137_9);
	INVX1 g_not_n1548 (n1548, not_n1548);
	BUFX2 g_n354 (and_not_pi014_2_pi054, n354);
	AND2X1 g_and_not_pi076_not_pi138_168070 (not_pi076, not_pi138_168070, and_not_pi076_not_pi138_168070);
	BUFX2 g_n1188 (and_pi026_pi053, n1188);
	INVX1 g_not_pi053_5 (pi053, not_pi053_5);
	AND2X1 g_and_n605_n607 (n607, n605, and_n605_n607);
	AND2X1 g_and_not_pi004_not_pi016 (not_pi004, not_pi016, and_not_pi004_not_pi016);
	BUFX2 g_n1504 (and_pi084_not_pi136_70, n1504);
	BUFX2 g_n559 (and_n449_n558, n559);
	BUFX2 g_n753 (and_not_pi058_not_n752, n753);
	INVX1 g_not_n1292 (n1292, not_n1292);
	BUFX2 g_n1048 (and_pi082_not_n1027, n1048);
	INVX1 g_not_n1084 (n1084, not_n1084);
	BUFX2 g_n1212 (and_not_pi053_8_n1211, n1212);
	AND2X1 g_and_not_pi110_6_n1419 (not_pi110_6, n1419, and_not_pi110_6_n1419);
	BUFX2 g_po060 (po060_driver, po060);
	AND2X1 g_and_not_pi043_not_pi047 (not_pi043, not_pi047, and_not_pi043_not_pi047);
	INVX1 g_not_n1297 (n1297, not_n1297);
	BUFX2 g_n1258 (and_not_n1255_not_n1257, n1258);
	INVX1 g_not_pi045_1 (pi045, not_pi045_1);
	INVX1 g_not_n992 (n992, not_n992);
	AND2X1 g_and_n640_n652 (n640, n652, and_n640_n652);
	BUFX2 g_n711 (and_not_n703_n710, n711);
	AND2X1 g_and_not_pi050_3_n404 (n404, not_pi050_3, and_not_pi050_3_n404);
	INVX1 g_not_n1603 (n1603, not_n1603);
	INVX1 g_not_n319 (n319, not_n319);
	AND2X1 g_and_not_pi110_2_n800 (n800, not_pi110_2, and_not_pi110_2_n800);
	BUFX2 g_n863 (and_not_n861_not_n862, n863);
	BUFX2 g_n660 (and_not_n648_n659, n660);
	INVX1 g_not_pi014_2 (pi014, not_pi014_2);
	BUFX2 g_n309 (and_not_pi056_n308, n309);
	AND2X1 g_and_not_pi053_2_not_pi058_1 (not_pi053_2, not_pi058_1, and_not_pi053_2_not_pi058_1);
	AND2X1 g_and_pi085_n787 (pi085, n787, and_pi085_n787);
	AND2X1 g_and_not_pi136_1_not_n1352 (not_pi136_1, not_n1352, and_not_pi136_1_not_n1352);
	INVX1 g_not_n690 (n690, not_n690);
	INVX1 g_not_pi096_0 (pi096, not_pi096_0);
	AND2X1 g_and_n502_n506 (n502, n506, and_n502_n506);
	BUFX2 g_n560 (and_n503_n559, n560);
	AND2X1 g_and_not_n1330_not_n1331 (not_n1330, not_n1331, and_not_n1330_not_n1331);
	AND2X1 g_and_not_n1338_not_n1339 (not_n1338, not_n1339, and_not_n1338_not_n1339);
	INVX1 g_not_pi048_1 (pi048, not_pi048_1);
	AND2X1 g_and_not_pi006_0_not_pi012_0 (not_pi012_0, not_pi006_0, and_not_pi006_0_not_pi012_0);
	BUFX2 g_n621 (and_pi016_pi054, n621);
	INVX1 g_not_pi143_0 (pi143, not_pi143_0);
	INVX1 g_not_pi136_8 (pi136, not_pi136_8);
	INVX1 g_not_pi106_6 (pi106, not_pi106_6);
	BUFX2 g_n1027 (and_n388_n391, n1027);
	AND2X1 g_and_not_n1448_not_n1449 (not_n1448, not_n1449, and_not_n1448_not_n1449);
	AND2X1 g_and_n487_n623 (n623, n487, and_n487_n623);
	AND2X1 g_and_pi026_n718 (n718, pi026, and_pi026_n718);
	OR2X1 g_or_pi129_n1314 (n1314, pi129, or_pi129_n1314);
	BUFX2 g_n442 (and_not_pi025_not_pi029, n442);
	BUFX2 g_n444 (and_n441_n443, n444);
	INVX1 g_not_n755 (n755, not_n755);
	INVX1 g_not_pi117 (pi117, not_pi117);
	BUFX2 g_n1141 (and_not_pi106_9_not_n943_0, n1141);
	AND2X1 g_and_not_n1290_not_n1292 (not_n1292, not_n1290, and_not_n1290_not_n1292);
	INVX1 g_not_pi002_0 (pi002, not_pi002_0);
	BUFX2 g_n1073 (and_n568_n572, n1073);
	INVX1 g_not_pi003_2326305139872070 (pi003, not_pi003_2326305139872070);
	INVX1 g_not_n733 (n733, not_n733);
	INVX1 g_not_n1549 (n1549, not_n1549);
	INVX1 g_not_pi008 (pi008, not_pi008);
	AND2X1 g_and_not_n353_not_n375 (not_n375, not_n353, and_not_n353_not_n375);
	BUFX2 g_n961 (and_n390_n960, n961);
	AND2X1 g_and_not_n829_not_n834 (not_n829, not_n834, and_not_n829_not_n834);
	AND2X1 g_and_not_n1255_not_n1257 (not_n1255, not_n1257, and_not_n1255_not_n1257);
	AND2X1 g_and_pi138_n1412 (pi138, n1412, and_pi138_n1412);
	INVX1 g_not_pi129_10045252112690790399992215344966975021805416861747224664747430 (pi129, not_pi129_10045252112690790399992215344966975021805416861747224664747430);
	INVX1 g_not_pi011_6 (pi011, not_pi011_6);
	BUFX2 g_n1132 (and_n934_n1131, n1132);
	AND2X1 g_and_not_pi106_4_not_n899 (not_pi106_4, not_n899, and_not_pi106_4_not_n899);
	INVX1 g_not_n873 (n873, not_n873);
	BUFX2 g_n464 (and_n445_n463, n464);
	BUFX2 g_n1094 (and_pi048_n1041, n1094);
	INVX1 g_not_pi026_9 (pi026, not_pi026_9);
	BUFX2 g_n1043 (and_n934_n1042, n1043);
	INVX1 g_not_n1541 (n1541, not_n1541);
	INVX1 g_not_pi129_302268019717750559482470516839540966128657419430 (pi129, not_pi129_302268019717750559482470516839540966128657419430);
	INVX1 g_not_pi136_7 (pi136, not_pi136_7);
	AND2X1 g_and_pi082_not_n927 (not_n927, pi082, and_pi082_not_n927);
	AND2X1 g_and_pi082_not_n919 (pi082, not_n919, and_pi082_not_n919);
	BUFX2 g_n1591 (and_not_n1589_not_n1590, n1591);
	AND2X1 g_and_n379_not_n1050 (n379, not_n1050, and_n379_not_n1050);
	INVX1 g_not_n1602 (n1602, not_n1602);
	AND2X1 g_and_n1606_n1607 (n1607, n1606, and_n1606_n1607);
	BUFX2 g_po115_driver (and_not_pi129_205005145156954906122290109080958673914396262484637238056070_not_n1446, po115_driver);
	BUFX2 g_n657 (and_pi082_not_n656, n657);
	AND2X1 g_and_pi045_n1041 (pi045, n1041, and_pi045_n1041);
	BUFX2 g_n1003 (and_n379_not_n1002, n1003);
	BUFX2 g_n1053 (and_not_pi046_2_not_n1052, n1053);
	BUFX2 g_po126_driver (and_not_pi129_492217353521848729599618551903381776068465426225614008572624070_n1586, po126_driver);
	INVX1 g_not_n1388 (n1388, not_n1388);
	BUFX2 g_n1283 (and_not_n1280_not_n1282, n1283);
	BUFX2 g_n1149 (and_not_pi053_5_not_n1148, n1149);
	BUFX2 g_po094 (po094_driver, po094);
	INVX1 g_not_pi052 (pi052, not_pi052);
	INVX1 g_not_pi048_2 (pi048, not_pi048_2);
	AND2X1 g_and_pi095_not_n1423 (not_n1423, pi095, and_pi095_not_n1423);
	AND2X1 g_and_pi137_not_n1463 (pi137, not_n1463, and_pi137_not_n1463);
	INVX1 g_not_n413 (n413, not_n413);
	AND2X1 g_and_not_pi048_3_not_n1084 (not_n1084, not_pi048_3, and_not_pi048_3_not_n1084);
	INVX1 g_not_n327 (n327, not_n327);
	AND2X1 g_and_not_pi028_n460 (not_pi028, n460, and_not_pi028_n460);
	BUFX2 g_n537 (and_pi018_n295, n537);
	BUFX2 g_n783 (and_pi027_n768, n783);
	AND2X1 g_and_not_pi026_6_not_pi100_1 (not_pi100_1, not_pi026_6, and_not_pi026_6_not_pi100_1);
	BUFX2 g_n857 (and_n838_n856, n857);
	BUFX2 g_n640 (and_n638_n639, n640);
	AND2X1 g_and_not_n379_2_not_n701 (not_n701, not_n379_2, and_not_n379_2_not_n701);
	INVX1 g_not_n770 (n770, not_n770);
	AND2X1 g_and_not_pi100_2_pi116 (pi116, not_pi100_2, and_not_pi100_2_pi116);
	AND2X1 g_and_pi082_not_n930 (pi082, not_n930, and_pi082_not_n930);
	BUFX2 g_n1580 (and_pi111_not_n1421_0, n1580);
	BUFX2 g_n1453 (and_pi093_pi138, n1453);
	INVX1 g_not_n950 (n950, not_n950);
	INVX1 g_not_n905 (n905, not_n905);
	INVX1 g_not_n1072 (n1072, not_n1072);
	AND2X1 g_and_not_n876_not_n877 (not_n877, not_n876, and_not_n876_not_n877);
	INVX1 g_not_n1214 (n1214, not_n1214);
	INVX1 g_not_n1361 (n1361, not_n1361);
	BUFX2 g_n1022 (and_not_n1020_not_n1021, n1022);
	BUFX2 g_n527 (and_not_pi010_2_pi022, n527);
	AND2X1 g_and_pi019_not_pi054_3430 (pi019, not_pi054_3430, and_pi019_not_pi054_3430);
	INVX1 g_not_pi096 (pi096, not_pi096);
	INVX1 g_not_n379_4 (n379, not_n379_4);
	INVX1 g_not_n1053 (n1053, not_n1053);
	AND2X1 g_and_pi037_n1360 (pi037, n1360, and_pi037_n1360);
	INVX1 g_not_n1540 (n1540, not_n1540);
	INVX1 g_not_n796_0 (n796, not_n796_0);
	BUFX2 g_n1218 (and_pi059_not_n1217, n1218);
	BUFX2 g_po078 (po078_driver, po078);
	INVX1 g_not_n898 (n898, not_n898);
	BUFX2 g_n918 (and_n406_n579, n918);
	BUFX2 g_n701 (and_pi082_not_n700, n701);
	AND2X1 g_and_not_pi017_1_pi054 (not_pi017_1, pi054, and_not_pi017_1_pi054);
	INVX1 g_not_pi044_2 (pi044, not_pi044_2);
	INVX1 g_not_n1048 (n1048, not_n1048);
	BUFX2 g_n1116 (and_not_n1114_not_n1115, n1116);
	AND2X1 g_and_n503_n525 (n525, n503, and_n503_n525);
	INVX1 g_not_n339 (n339, not_n339);
	AND2X1 g_and_not_pi053_8_n1211 (n1211, not_pi053_8, and_not_pi053_8_n1211);
	AND2X1 g_and_pi087_not_pi138_3 (pi087, not_pi138_3, and_pi087_not_pi138_3);
	AND2X1 g_and_not_pi003_19773267430_n1153 (not_pi003_19773267430, n1153, and_not_pi003_19773267430_n1153);
	BUFX2 g_po092 (po092_driver, po092);
	INVX1 g_not_n314 (n314, not_n314);
	BUFX2 g_n1407 (and_pi093_not_n1386_4, n1407);
	INVX1 g_not_pi050_3 (pi050, not_pi050_3);
	INVX1 g_not_pi129_8 (pi129, not_pi129_8);
	AND2X1 g_and_n1251_n1324 (n1251, n1324, and_n1251_n1324);
	BUFX2 g_po042_driver (and_n786_n788, po042_driver);
	AND2X1 g_and_not_pi116_0_n747 (not_pi116_0, n747, and_not_pi116_0_n747);
	BUFX2 g_n1158 (and_pi082_not_n1157, n1158);
	OR2X1 g_or_pi129_n1258 (pi129, n1258, or_pi129_n1258);
	INVX1 g_not_n975 (n975, not_n975);
	INVX1 g_not_n379_70 (n379, not_n379_70);
	BUFX2 g_n1379 (and_not_n1377_not_n1378, n1379);
	BUFX2 g_po018 (po018_driver, po018);
	INVX1 g_not_pi096_2 (pi096, not_pi096_2);
	AND2X1 g_and_not_n740_not_n741 (not_n740, not_n741, and_not_n740_not_n741);
	INVX1 g_not_n1183 (n1183, not_n1183);
	AND2X1 g_and_not_n1511_not_n1512 (not_n1511, not_n1512, and_not_n1511_not_n1512);
	BUFX2 g_po091 (po091_driver, po091);
	AND2X1 g_and_pi026_not_pi027_5 (not_pi027_5, pi026, and_pi026_not_pi027_5);
	AND2X1 g_and_n638_n954 (n954, n638, and_n638_n954);
	INVX1 g_not_n379 (n379, not_n379);
	INVX1 g_not_n1474 (n1474, not_n1474);
	INVX1 g_not_n1174 (n1174, not_n1174);
	AND2X1 g_and_not_pi129_13410686196639649008070_not_n908 (not_pi129_13410686196639649008070, not_n908, and_not_pi129_13410686196639649008070_not_n908);
	INVX1 g_not_n987 (n987, not_n987);
	BUFX2 g_n653 (and_n640_n652, n653);
	BUFX2 g_n1137 (and_not_n940_not_n1136, n1137);
	AND2X1 g_and_pi057_not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490 (pi057, not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490, and_pi057_not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490);
	INVX1 g_not_n806 (n806, not_n806);
	INVX1 g_not_pi000 (pi000, not_pi000);
	AND2X1 g_and_n357_n549 (n549, n357, and_n357_n549);
	AND2X1 g_and_pi026_not_pi058_6 (not_pi058_6, pi026, and_pi026_not_pi058_6);
	INVX1 g_not_n635 (n635, not_n635);
	BUFX2 g_n1524 (and_not_pi136_3430_not_n1523, n1524);
	AND2X1 g_and_not_n790_not_n791 (not_n790, not_n791, and_not_n790_not_n791);
	BUFX2 g_n665 (and_pi019_n664, n665);
	AND2X1 g_and_not_pi058_7_n1175 (not_pi058_7, n1175, and_not_pi058_7_n1175);
	BUFX2 g_n1549 (and_not_n1544_not_n1548, n1549);
	AND2X1 g_and_n776_n801 (n776, n801, and_n776_n801);
	AND2X1 g_and_not_pi129_2115876138024253916377293617876786762900601936010_not_n1383 (not_pi129_2115876138024253916377293617876786762900601936010, not_n1383, and_not_pi129_2115876138024253916377293617876786762900601936010_not_n1383);
	INVX1 g_not_pi054_1176490 (pi054, not_pi054_1176490);
	INVX1 g_not_pi016_1 (pi016, not_pi016_1);
	AND2X1 g_and_not_pi044_2_n649 (not_pi044_2, n649, and_not_pi044_2_n649);
	INVX1 g_not_n1282 (n1282, not_n1282);
	AND2X1 g_and_n344_n348 (n344, n348, and_n344_n348);
	BUFX2 g_po014_driver (pi128, po014_driver);
	BUFX2 g_po010 (po010_driver, po010);
	BUFX2 g_n505 (and_n448_n504, n505);
	BUFX2 g_n1008 (and_pi082_not_n1007, n1008);
	AND2X1 g_and_pi049_n411 (n411, pi049, and_pi049_n411);
	AND2X1 g_and_n314_n322 (n314, n322, and_n314_n322);
	BUFX2 g_n387 (and_not_pi041_not_pi046, n387);
	INVX1 g_not_pi005_5 (pi005, not_pi005_5);
	INVX1 g_not_n834 (n834, not_n834);
	BUFX2 g_po095_driver (and_not_pi129_17984650426474121466202803405696493492512490_not_n1336, po095_driver);
	BUFX2 g_n1198 (and_not_n1195_not_n1197, n1198);
	BUFX2 g_n1001 (and_n385_n698, n1001);
	BUFX2 g_po012 (po012_driver, po012);
	INVX1 g_not_n668 (n668, not_n668);
	BUFX2 g_n482 (and_n478_n481, n482);
	BUFX2 g_n1097 (and_not_pi129_185621159210175743024531636712070_not_n1096, n1097);
	BUFX2 g_n1344 (and_not_n1342_not_n1343, n1344);
	INVX1 g_not_pi129_47475615099430 (pi129, not_pi129_47475615099430);
	AND2X1 g_and_not_pi004_1_not_pi018_3 (not_pi004_1, not_pi018_3, and_not_pi004_1_not_pi018_3);
	INVX1 g_not_n1486 (n1486, not_n1486);
	BUFX2 g_po013_driver (pi130, po013_driver);
	BUFX2 g_n1560 (and_not_n1555_not_n1559, n1560);
	INVX1 g_not_pi024_1 (pi024, not_pi024_1);
	BUFX2 g_n920 (and_n918_n919, n920);
	AND2X1 g_and_not_pi129_5585458640832840070_not_n880 (not_pi129_5585458640832840070, not_n880, and_not_pi129_5585458640832840070_not_n880);
	INVX1 g_not_pi129_32199057558131797268376070 (pi129, not_pi129_32199057558131797268376070);
	AND2X1 g_and_n332_n500 (n332, n500, and_n332_n500);
	INVX1 g_not_n1226 (n1226, not_n1226);
	INVX1 g_not_pi007_3 (pi007, not_pi007_3);
	BUFX2 g_n1584 (and_n1581_n1583, n1584);
	BUFX2 g_n1272 (and_pi066_not_n1271, n1272);
	BUFX2 g_po000_driver (pi108, po000_driver);
	BUFX2 g_n1112 (and_n380_n1111, n1112);
	AND2X1 g_and_pi146_n1386 (pi146, n1386, and_pi146_n1386);
	INVX1 g_not_n1449 (n1449, not_n1449);
	INVX1 g_not_n765 (n765, not_n765);
	AND2X1 g_and_pi082_not_n1325_3 (not_n1325_3, pi082, and_pi082_not_n1325_3);
	BUFX2 g_n1069 (and_n408_n927, n1069);
	AND2X1 g_and_pi082_not_n575 (not_n575, pi082, and_pi082_not_n575);
	INVX1 g_not_n1616 (n1616, not_n1616);
	AND2X1 g_and_pi082_not_n1113 (not_n1113, pi082, and_pi082_not_n1113);
	BUFX2 g_n734 (and_not_n721_not_n733, n734);
	BUFX2 g_n799 (and_pi028_not_n798, n799);
	INVX1 g_not_pi049_1 (pi049, not_pi049_1);
	AND2X1 g_and_pi082_not_n1121 (pi082, not_n1121, and_pi082_not_n1121);
	BUFX2 g_n739 (and_not_n718_not_n738, n739);
	BUFX2 g_n727 (and_pi025_not_n726, n727);
	BUFX2 g_n834 (and_n724_not_n833, n834);
	AND2X1 g_and_not_pi005_5_n596 (not_pi005_5, n596, and_not_pi005_5_n596);
	AND2X1 g_and_n401_n926 (n926, n401, and_n401_n926);
	INVX1 g_not_n1506 (n1506, not_n1506);
	BUFX2 g_n345 (and_not_pi007_2_not_pi013_2, n345);
	AND2X1 g_and_not_n1312_not_n1313 (not_n1312, not_n1313, and_not_n1312_not_n1313);
	AND2X1 g_and_not_pi026_0_not_pi085_1 (not_pi026_0, not_pi085_1, and_not_pi026_0_not_pi085_1);
	INVX1 g_not_pi129_273687473400809163430 (pi129, not_pi129_273687473400809163430);
	INVX1 g_not_pi072 (pi072, not_pi072);
	BUFX2 g_n1566 (and_pi030_n1360, n1566);
	BUFX2 g_n866 (and_not_n864_not_n865, n866);
	AND2X1 g_and_not_pi085_not_pi110 (not_pi110, not_pi085, and_not_pi085_not_pi110);
	AND2X1 g_and_not_n864_not_n865 (not_n865, not_n864, and_not_n864_not_n865);
	OR2X1 g_or_pi129_n1318 (n1318, pi129, or_pi129_n1318);
	BUFX2 g_n962 (and_not_pi129_32199057558131797268376070_not_n961, n962);
	AND2X1 g_and_n390_n977 (n390, n977, and_n390_n977);
	BUFX2 g_n360 (and_pi006_pi012, n360);
	OR2X1 g_or_pi129_n1288 (pi129, n1288, or_pi129_n1288);
	BUFX2 g_n476 (and_not_pi007_6_n449, n476);
	AND2X1 g_and_not_n362_not_n363 (not_n362, not_n363, and_not_n362_not_n363);
	AND2X1 g_and_n293_n296 (n293, n296, and_n293_n296);
	BUFX2 g_n932 (and_not_n379_3_not_n931, n932);
	AND2X1 g_and_not_n1300_not_n1301 (not_n1300, not_n1301, and_not_n1300_not_n1301);
	INVX1 g_not_n370 (n370, not_n370);
	INVX1 g_not_n1038 (n1038, not_n1038);
	AND2X1 g_and_not_n726_1_n787 (not_n726_1, n787, and_not_n726_1_n787);
	BUFX2 g_n1274 (and_not_n1272_not_n1273, n1274);
	BUFX2 g_n1206 (and_pi116_not_n796_0, n1206);
	BUFX2 g_po100 (po100_driver, po100);
	BUFX2 g_n325 (and_not_pi010_not_n324, n325);
	BUFX2 g_n393 (and_n389_n392, n393);
	AND2X1 g_and_not_pi058_8_not_n1190 (not_pi058_8, not_n1190, and_not_pi058_8_not_n1190);
	BUFX2 g_n1028 (and_n1026_n1027, n1028);
	AND2X1 g_and_not_pi026_168070_n1375 (not_pi026_168070, n1375, and_not_pi026_168070_n1375);
	INVX1 g_not_n1473 (n1473, not_n1473);
	INVX1 g_not_pi013_1 (pi013, not_pi013_1);
	BUFX2 g_n297 (and_n293_n296, n297);
	INVX1 g_not_pi109_3 (pi109, not_pi109_3);
	BUFX2 g_n1127 (and_n927_n1126, n1127);
	INVX1 g_not_pi026_24010 (pi026, not_pi026_24010);
	AND2X1 g_and_not_n582_not_n588 (not_n588, not_n582, and_not_n582_not_n588);
	BUFX2 g_po076_driver (and_not_pi129_52433383167563036344614587188619514555430_n1241, po076_driver);
	AND2X1 g_and_not_pi129_52433383167563036344614587188619514555430_n1241 (not_pi129_52433383167563036344614587188619514555430, n1241, and_not_pi129_52433383167563036344614587188619514555430_n1241);
	BUFX2 g_n1397 (and_not_n1395_not_n1396, n1397);
	INVX1 g_not_n1092 (n1092, not_n1092);
	BUFX2 g_n691 (and_pi082_not_n690, n691);
	AND2X1 g_and_not_pi129_0_not_n376 (not_pi129_0, not_n376, and_not_pi129_0_not_n376);
	AND2X1 g_and_not_pi129_8235430_not_n625 (not_n625, not_pi129_8235430, and_not_pi129_8235430_not_n625);
	BUFX2 g_n1004 (and_not_n1000_not_n1003, n1004);
	INVX1 g_not_pi129_2 (pi129, not_pi129_2);
	INVX1 g_not_pi054_6 (pi054, not_pi054_6);
	INVX1 g_not_n584 (n584, not_n584);
	AND2X1 g_and_pi046_pi082 (pi046, pi082, and_pi046_pi082);
	BUFX2 g_n1306 (and_not_n1304_not_n1305, n1306);
	AND2X1 g_and_n408_n699 (n699, n408, and_n408_n699);
	INVX1 g_not_pi136_9 (pi136, not_pi136_9);
	BUFX2 g_n991 (and_n638_n990, n991);
	INVX1 g_not_n731 (n731, not_n731);
	INVX1 g_not_n882 (n882, not_n882);
	AND2X1 g_and_pi042_n934 (n934, pi042, and_pi042_n934);
	BUFX2 g_po015 (po015_driver, po015);
	AND2X1 g_and_not_n1020_not_n1021 (not_n1020, not_n1021, and_not_n1020_not_n1021);
	INVX1 g_not_pi129_24118650322570587750381309043265707027354805885055086420058579430 (pi129, not_pi129_24118650322570587750381309043265707027354805885055086420058579430);
	BUFX2 g_po122_driver (or_n1543_n1550, po122_driver);
	BUFX2 g_po030_driver (and_not_pi129_24010_not_n593, po030_driver);
	INVX1 g_not_pi018_0 (pi018, not_pi018_0);
	INVX1 g_not_pi129_138412872010 (pi129, not_pi129_138412872010);
	AND2X1 g_and_not_pi110_7_not_pi120 (not_pi120, not_pi110_7, and_not_pi110_7_not_pi120);
	BUFX2 g_n1136 (and_pi051_not_pi109_7, n1136);
	INVX1 g_not_n1565 (n1565, not_n1565);
	INVX1 g_not_pi047_0 (pi047, not_pi047_0);
	INVX1 g_not_pi014_0 (pi014, not_pi014_0);
	INVX1 g_not_pi129_445676403263631959001900459745680070 (pi129, not_pi129_445676403263631959001900459745680070);
	AND2X1 g_and_not_n1459_not_n1460 (not_n1460, not_n1459, and_not_n1459_not_n1460);
	INVX1 g_not_pi002_3 (pi002, not_pi002_3);
	BUFX2 g_n1002 (and_pi082_not_n1001, n1002);
	INVX1 g_not_pi003_5585458640832840070 (pi003, not_pi003_5585458640832840070);
	INVX1 g_not_pi054_2 (pi054, not_pi054_2);
	AND2X1 g_and_pi010_n291 (pi010, n291, and_pi010_n291);
	BUFX2 g_n397 (and_not_pi065_n396, n397);
	INVX1 g_not_n1295 (n1295, not_n1295);
	AND2X1 g_and_not_n1068_n1078 (n1078, not_n1068, and_not_n1068_n1078);
	BUFX2 g_n719 (and_pi085_n718, n719);
	AND2X1 g_and_not_n1489_not_n1490 (not_n1489, not_n1490, and_not_n1489_not_n1490);
	BUFX2 g_n1383 (and_not_n1381_not_n1382, n1383);
	AND2X1 g_and_not_n767_not_n769 (not_n767, not_n769, and_not_n767_not_n769);
	BUFX2 g_n699 (and_n401_n698, n699);
	AND2X1 g_and_pi111_pi138 (pi111, pi138, and_pi111_pi138);
	INVX1 g_not_pi053_6 (pi053, not_pi053_6);
	BUFX2 g_n512 (and_not_pi010_1_n449, n512);
	INVX1 g_not_n1117 (n1117, not_n1117);
	INVX1 g_not_n404 (n404, not_n404);
	AND2X1 g_and_not_pi085_4_not_n738_0 (not_pi085_4, not_n738_0, and_not_pi085_4_not_n738_0);
	INVX1 g_not_n379_8 (n379, not_n379_8);
	AND2X1 g_and_not_pi005_1_n332 (not_pi005_1, n332, and_not_pi005_1_n332);
	BUFX2 g_n404 (and_n390_n403, n404);
	INVX1 g_not_n1132 (n1132, not_n1132);
	INVX1 g_not_n1437 (n1437, not_n1437);
	INVX1 g_not_pi003_332329305696010 (pi003, not_pi003_332329305696010);
	INVX1 g_not_n1536 (n1536, not_n1536);
	AND2X1 g_and_n316_n318 (n316, n318, and_n316_n318);
	INVX1 g_not_pi012_2 (pi012, not_pi012_2);
	BUFX2 g_n1089 (and_n408_n1088, n1089);
	INVX1 g_not_pi003_1 (pi003, not_pi003_1);
	INVX1 g_not_pi085_4 (pi085, not_pi085_4);
	INVX1 g_not_n1003 (n1003, not_n1003);
	INVX1 g_not_pi043_2 (pi043, not_pi043_2);
	INVX1 g_not_pi007_1 (pi007, not_pi007_1);
	INVX1 g_not_n823 (n823, not_n823);
	BUFX2 g_n893 (and_not_pi106_3_not_n892, n893);
	AND2X1 g_and_not_n1023_n1024 (n1024, not_n1023, and_not_n1023_n1024);
	AND2X1 g_and_pi097_not_pi110_3 (not_pi110_3, pi097, and_pi097_not_pi110_3);
	INVX1 g_not_pi122_1 (pi122, not_pi122_1);
	AND2X1 g_and_n1583_n1600 (n1600, n1583, and_n1583_n1600);
	BUFX2 g_po052_driver (and_not_pi129_93874803376477543056490_not_n915, po052_driver);
	BUFX2 g_po099 (po099_driver, po099);
	BUFX2 g_po053 (po053_driver, po053);
	INVX1 g_not_n1351 (n1351, not_n1351);
	AND2X1 g_and_pi088_not_n1386 (pi088, not_n1386, and_pi088_not_n1386);
	AND2X1 g_and_n786_n788 (n788, n786, and_n786_n788);
	BUFX2 g_n536 (and_n448_n535, n536);
	BUFX2 g_n986 (and_pi082_not_n985, n986);
	BUFX2 g_po049 (po049_driver, po049);
	INVX1 g_not_pi026_0 (pi026, not_pi026_0);
	INVX1 g_not_n746 (n746, not_n746);
	INVX1 g_not_pi013_5 (pi013, not_pi013_5);
	INVX1 g_not_n376 (n376, not_n376);
	INVX1 g_not_n1055 (n1055, not_n1055);
	AND2X1 g_and_not_pi082_n379 (n379, not_pi082, and_not_pi082_n379);
	INVX1 g_not_n1190 (n1190, not_n1190);
	BUFX2 g_n1357 (and_pi087_not_pi138_3, n1357);
	BUFX2 g_po002_driver (pi104, po002_driver);
	AND2X1 g_and_pi099_not_n1386_6 (not_n1386_6, pi099, and_pi099_not_n1386_6);
	BUFX2 g_n618 (and_not_pi129_1176490_not_n617, n618);
	INVX1 g_not_n1456 (n1456, not_n1456);
	BUFX2 g_n1577 (and_not_pi129_70316764788835532799945507414768825152637918032230572653232010_not_n1576, n1577);
	AND2X1 g_and_n408_n585 (n408, n585, and_n408_n585);
	INVX1 g_not_pi115_0 (pi115, not_pi115_0);
	OR2X1 g_or_n1561_n1568 (n1561, n1568, or_n1561_n1568);
	INVX1 g_not_n996 (n996, not_n996);
	INVX1 g_not_n1386_1 (n1386, not_n1386_1);
	AND2X1 g_and_not_n1108_not_n1112 (not_n1112, not_n1108, and_not_n1108_not_n1112);
	AND2X1 g_and_pi030_pi109 (pi030, pi109, and_pi030_pi109);
	AND2X1 g_and_not_pi007_4_n332 (not_pi007_4, n332, and_not_pi007_4_n332);
	BUFX2 g_n1185 (and_not_pi129_21838143759917965991093122527538323430_not_n1184, n1185);
	INVX1 g_not_n364 (n364, not_n364);
	AND2X1 g_and_n675_n680 (n675, n680, and_n675_n680);
	BUFX2 g_n1110 (and_n1100_not_n1109, n1110);
	AND2X1 g_and_not_n1169_not_n1171 (not_n1171, not_n1169, and_not_n1169_not_n1171);
	BUFX2 g_n981 (and_not_n975_n980, n981);
	INVX1 g_not_n1325_4 (n1325, not_n1325_4);
	INVX1 g_not_pi012_6 (pi012, not_pi012_6);
	AND2X1 g_and_not_n662_not_n668 (not_n668, not_n662, and_not_n662_not_n668);
	INVX1 g_not_n1570 (n1570, not_n1570);
	AND2X1 g_and_not_n823_not_n825 (not_n823, not_n825, and_not_n823_not_n825);
	AND2X1 g_and_not_n1350_not_n1351 (not_n1351, not_n1350, and_not_n1350_not_n1351);
	BUFX2 g_n435 (and_n432_n434, n435);
	BUFX2 g_n1211 (and_not_pi003_6782230728490_n1210, n1211);
	AND2X1 g_and_n927_n1017 (n927, n1017, and_n927_n1017);
	BUFX2 g_n1483 (and_not_n1481_not_n1482, n1483);
	INVX1 g_not_pi129_52433383167563036344614587188619514555430 (pi129, not_pi129_52433383167563036344614587188619514555430);
	OR2X1 g_or_n1543_n1550 (n1550, n1543, or_n1543_n1550);
	INVX1 g_not_pi113 (pi113, not_pi113);
	BUFX2 g_n507 (and_n502_n506, n507);
	BUFX2 g_n1430 (and_not_n1428_not_n1429, n1430);
	INVX1 g_not_n628 (n628, not_n628);
	INVX1 g_not_n1051 (n1051, not_n1051);
	INVX1 g_not_n1401 (n1401, not_n1401);
	INVX1 g_not_n1421_0 (n1421, not_n1421_0);
	AND2X1 g_and_pi034_not_pi109_3 (not_pi109_3, pi034, and_pi034_not_pi109_3);
	INVX1 g_not_n1493 (n1493, not_n1493);
	INVX1 g_not_pi026_5 (pi026, not_pi026_5);
	BUFX2 g_po039 (po039_driver, po039);
	BUFX2 g_n601 (and_not_n595_not_n600, n601);
	BUFX2 g_n707 (and_n390_n706, n707);
	BUFX2 g_n1312 (and_pi075_not_n1271_4, n1312);
	AND2X1 g_and_pi076_n974 (n974, pi076, and_pi076_n974);
	AND2X1 g_and_pi136_not_n1454 (not_n1454, pi136, and_pi136_not_n1454);
	BUFX2 g_n376 (and_not_n353_not_n375, n376);
	BUFX2 g_n1131 (and_pi050_n1041, n1131);
	BUFX2 g_n1543 (and_not_pi137_9_not_n1542, n1543);
	INVX1 g_not_pi047_1 (pi047, not_pi047_1);
	INVX1 g_not_n1178 (n1178, not_n1178);
	AND2X1 g_and_not_n1432_not_n1433 (not_n1433, not_n1432, and_not_n1432_not_n1433);
	INVX1 g_not_pi048_0 (pi048, not_pi048_0);
	INVX1 g_not_pi051_1 (pi051, not_pi051_1);
	AND2X1 g_and_n390_n650 (n390, n650, and_n390_n650);
	BUFX2 g_po120_driver (or_n1520_n1527, po120_driver);
	AND2X1 g_and_not_pi040_1_not_pi042_0 (not_pi042_0, not_pi040_1, and_not_pi040_1_not_pi042_0);
	AND2X1 g_and_not_n703_n710 (n710, not_n703, and_not_n703_n710);
	AND2X1 g_and_n1251_n1385 (n1251, n1385, and_n1251_n1385);
	BUFX2 g_po108 (po108_driver, po108);
	INVX1 g_not_n940_0 (n940, not_n940_0);
	BUFX2 g_n1396 (and_pi142_n1386, n1396);
	BUFX2 g_n508 (and_not_n498_not_n507, n508);
	AND2X1 g_and_pi087_not_n1325_6 (pi087, not_n1325_6, and_pi087_not_n1325_6);
	INVX1 g_not_n1221 (n1221, not_n1221);
	INVX1 g_not_n1194 (n1194, not_n1194);
	AND2X1 g_and_pi091_n1249 (n1249, pi091, and_pi091_n1249);
	INVX1 g_not_pi082 (pi082, not_pi082);
	BUFX2 g_n514 (and_n503_n513, n514);
	AND2X1 g_and_not_pi059_n356 (n356, not_pi059, and_not_pi059_n356);
	AND2X1 g_and_pi078_not_pi136_8 (not_pi136_8, pi078, and_pi078_not_pi136_8);
	BUFX2 g_n901 (and_not_n896_not_n900, n901);
	AND2X1 g_and_pi131_n1245 (n1245, pi131, and_pi131_n1245);
	AND2X1 g_and_n927_n971 (n971, n927, and_n927_n971);
	INVX1 g_not_pi063 (pi063, not_pi063);
	BUFX2 g_n1607 (and_not_pi007_10_not_pi009_6, n1607);
	INVX1 g_not_pi116_70 (pi116, not_pi116_70);
	BUFX2 g_n1538 (and_not_pi076_not_pi138_168070, n1538);
	AND2X1 g_and_pi089_pi106 (pi089, pi106, and_pi089_pi106);
	AND2X1 g_and_not_n953_n963 (n963, not_n953, and_not_n953_n963);
	AND2X1 g_and_not_pi106_8_n1137 (n1137, not_pi106_8, and_not_pi106_8_n1137);
	AND2X1 g_and_not_n810_not_n811 (not_n810, not_n811, and_not_n810_not_n811);
	BUFX2 g_n1424 (and_pi095_not_n1423, n1424);
	INVX1 g_not_n1257 (n1257, not_n1257);
	AND2X1 g_and_not_n1452_not_n1453 (not_n1453, not_n1452, and_not_n1452_not_n1453);
	BUFX2 g_n1494 (and_not_pi138_9_not_n1493, n1494);
	AND2X1 g_and_not_pi016_0_pi054 (not_pi016_0, pi054, and_not_pi016_0_pi054);
	BUFX2 g_n1278 (and_not_n1276_not_n1277, n1278);
	BUFX2 g_po136_driver (and_not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070_n1623, po136_driver);
	BUFX2 g_po077 (po077_driver, po077);
	INVX1 g_not_n1122 (n1122, not_n1122);
	BUFX2 g_n1562 (and_pi086_not_pi138_403536070, n1562);
	BUFX2 g_n1066 (and_n379_not_n1065, n1066);
	AND2X1 g_and_pi146_n1325 (pi146, n1325, and_pi146_n1325);
	BUFX2 g_n612 (and_not_pi011_5_n311, n612);
	BUFX2 g_n1184 (and_not_n1181_not_n1183, n1184);
	INVX1 g_not_n1157 (n1157, not_n1157);
	INVX1 g_not_pi003_797922662976120010 (pi003, not_pi003_797922662976120010);
	BUFX2 g_po044_driver (and_not_pi003_2824752490_n859, po044_driver);
	AND2X1 g_and_not_n742_n743 (n743, not_n742, and_not_n742_n743);
	INVX1 g_not_pi129_5585458640832840070 (pi129, not_pi129_5585458640832840070);
	BUFX2 g_n668 (and_n487_n667, n668);
	BUFX2 g_n347 (and_n345_n346, n347);
	INVX1 g_not_pi040_0 (pi040, not_pi040_0);
	AND2X1 g_and_pi082_not_n407 (not_n407, pi082, and_pi082_not_n407);
	INVX1 g_not_n1148 (n1148, not_n1148);
	INVX1 g_not_n1591 (n1591, not_n1591);
	INVX1 g_not_pi059_0 (pi059, not_pi059_0);
	INVX1 g_not_pi138_0 (pi138, not_pi138_0);
	BUFX2 g_n333 (and_n331_n332, n333);
	BUFX2 g_n678 (and_pi005_not_pi007_9, n678);
	BUFX2 g_po011 (po011_driver, po011);
	INVX1 g_not_pi058_5 (pi058, not_pi058_5);
	INVX1 g_not_n337 (n337, not_n337);
	INVX1 g_not_pi052_0 (pi052, not_pi052_0);
	INVX1 g_not_n1271_3 (n1271, not_n1271_3);
	INVX1 g_not_n1560 (n1560, not_n1560);
	BUFX2 g_n1322 (and_not_n1320_not_n1321, n1322);
	INVX1 g_not_n1483 (n1483, not_n1483);
	AND2X1 g_and_not_pi027_0_n749 (n749, not_pi027_0, and_not_pi027_0_n749);
	BUFX2 g_n1246 (and_pi131_n1245, n1246);
	INVX1 g_not_n1356 (n1356, not_n1356);
	AND2X1 g_and_not_pi008_1_not_pi011_1 (not_pi011_1, not_pi008_1, and_not_pi008_1_not_pi011_1);
	INVX1 g_not_pi106_5 (pi106, not_pi106_5);
	BUFX2 g_po137_driver (or_pi129_pi134, po137_driver);
	AND2X1 g_and_pi082_not_pi138_7 (pi082, not_pi138_7, and_pi082_not_pi138_7);
	BUFX2 g_n956 (and_n927_n955, n956);
	INVX1 g_not_n317 (n317, not_n317);
	INVX1 g_not_n728_0 (n728, not_n728_0);
	BUFX2 g_n1174 (and_not_pi053_6_not_n1173, n1174);
	AND2X1 g_and_not_pi003_1915812313805664144010_not_n1628 (not_n1628, not_pi003_1915812313805664144010, and_not_pi003_1915812313805664144010_not_n1628);
	AND2X1 g_and_not_n1048_not_n1051 (not_n1051, not_n1048, and_not_n1048_not_n1051);
	INVX1 g_not_pi129_1 (pi129, not_pi129_1);
	BUFX2 g_po028 (po028_driver, po028);
	INVX1 g_not_n1462 (n1462, not_n1462);
	AND2X1 g_and_pi116_n1573 (pi116, n1573, and_pi116_n1573);
	INVX1 g_not_n802 (n802, not_n802);
	INVX1 g_not_n1172 (n1172, not_n1172);
	AND2X1 g_and_not_n1248_not_n1252 (not_n1252, not_n1248, and_not_n1248_not_n1252);
	INVX1 g_not_n1231 (n1231, not_n1231);
	AND2X1 g_and_pi136_n1243 (n1243, pi136, and_pi136_n1243);
	INVX1 g_not_n1408 (n1408, not_n1408);
	AND2X1 g_and_not_pi003_39098210485829880490_n1609 (n1609, not_pi003_39098210485829880490, and_not_pi003_39098210485829880490_n1609);
	BUFX2 g_n948 (and_n579_n919, n948);
	AND2X1 g_and_not_pi003_70_n618 (n618, not_pi003_70, and_not_pi003_70_n618);
	BUFX2 g_po064_driver (and_not_pi129_1299348114471230201171721456984490_not_n1117, po064_driver);
	AND2X1 g_and_pi090_pi106 (pi090, pi106, and_pi090_pi106);
	BUFX2 g_n1115 (and_pi049_n411, n1115);
	AND2X1 g_and_pi082_not_n656 (pi082, not_n656, and_pi082_not_n656);
	AND2X1 g_and_not_n1481_not_n1482 (not_n1482, not_n1481, and_not_n1481_not_n1482);
	BUFX2 g_po002 (po002_driver, po002);
	AND2X1 g_and_not_pi025_not_pi029 (not_pi029, not_pi025, and_not_pi025_not_pi029);
	BUFX2 g_n919 (and_n385_n697, n919);
	INVX1 g_not_pi129_13410686196639649008070 (pi129, not_pi129_13410686196639649008070);
	BUFX2 g_n771 (and_not_pi129_47475615099430_not_n770, n771);
	AND2X1 g_and_not_n1496_not_n1497 (not_n1496, not_n1497, and_not_n1496_not_n1497);
	BUFX2 g_n710 (and_not_pi129_968890104070_not_n709, n710);
	BUFX2 g_n406 (and_not_pi041_0_n405, n406);
	AND2X1 g_and_not_pi054_1176490_not_pi113_0 (not_pi054_1176490, not_pi113_0, and_not_pi054_1176490_not_pi113_0);
	AND2X1 g_and_not_pi002_4_not_pi047_4 (not_pi047_4, not_pi002_4, and_not_pi002_4_not_pi047_4);
	AND2X1 g_and_not_pi117_not_pi122_0 (not_pi122_0, not_pi117, and_not_pi117_not_pi122_0);
	INVX1 g_not_n1246 (n1246, not_n1246);
	AND2X1 g_and_not_pi004_2_not_pi012_6 (not_pi004_2, not_pi012_6, and_not_pi004_2_not_pi012_6);
	BUFX2 g_n540 (and_n538_n539, n540);
	BUFX2 g_n319 (and_n316_n318, n319);
	BUFX2 g_n1392 (and_pi140_n1386, n1392);
	INVX1 g_not_pi026_10 (pi026, not_pi026_10);
	INVX1 g_not_n377 (n377, not_n377);
	BUFX2 g_n728 (and_pi026_pi116, n728);
	BUFX2 g_po032 (po032_driver, po032);
	BUFX2 g_po081_driver (or_pi129_n1274, po081_driver);
	BUFX2 g_n466 (and_n448_n465, n466);
	BUFX2 g_po103 (po103_driver, po103);
	AND2X1 g_and_n291_n292 (n292, n291, and_n291_n292);
	BUFX2 g_n310 (and_not_pi056_0_not_n301, n310);
	BUFX2 g_n652 (and_n649_n651, n652);
	AND2X1 g_and_pi008_pi021 (pi021, pi008, and_pi008_pi021);
	AND2X1 g_and_n311_n341 (n311, n341, and_n311_n341);
	BUFX2 g_n825 (and_n819_n824, n825);
	BUFX2 g_n934 (and_not_pi044_1_pi082, n934);
	AND2X1 g_and_n1026_n1027 (n1027, n1026, and_n1026_n1027);
	INVX1 g_not_pi003_19773267430 (pi003, not_pi003_19773267430);
	INVX1 g_not_n1273 (n1273, not_n1273);
	INVX1 g_not_n890 (n890, not_n890);
	AND2X1 g_and_pi138_n1246 (n1246, pi138, and_pi138_n1246);
	BUFX2 g_n1445 (and_pi144_n1414, n1445);
	AND2X1 g_and_not_pi026_not_n720 (not_pi026, not_n720, and_not_pi026_not_n720);
	AND2X1 g_and_not_pi136_1176490_not_n1558 (not_n1558, not_pi136_1176490, and_not_pi136_1176490_not_n1558);
	BUFX2 g_n968 (and_not_n965_not_n967, n968);
	AND2X1 g_and_pi006_pi012 (pi006, pi012, and_pi006_pi012);
	AND2X1 g_and_pi064_not_n1247_1 (pi064, not_n1247_1, and_pi064_not_n1247_1);
	INVX1 g_not_n717 (n717, not_n717);
	INVX1 g_not_n1104 (n1104, not_n1104);
	AND2X1 g_and_not_pi115_0_not_n1421_2 (not_pi115_0, not_n1421_2, and_not_pi115_0_not_n1421_2);
	INVX1 g_not_n1386 (n1386, not_n1386);
	AND2X1 g_and_not_pi058_2_not_n822 (not_n822, not_pi058_2, and_not_pi058_2_not_n822);
	AND2X1 g_and_not_n648_n659 (n659, not_n648, and_not_n648_n659);
	INVX1 g_not_n1227 (n1227, not_n1227);
	BUFX2 g_po033_driver (and_not_pi003_490_n626, po033_driver);
	BUFX2 g_po026 (po026_driver, po026);
	BUFX2 g_n1119 (and_pi082_not_n404, n1119);
	BUFX2 g_n957 (and_pi082_not_n956, n957);
	INVX1 g_not_n1334 (n1334, not_n1334);
	AND2X1 g_and_not_n1356_not_n1357 (not_n1356, not_n1357, and_not_n1356_not_n1357);
	AND2X1 g_and_not_pi053_4_not_n841 (not_n841, not_pi053_4, and_not_pi053_4_not_n841);
	INVX1 g_not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070 (pi129, not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070);
	BUFX2 g_po130 (po130_driver, po130);
	AND2X1 g_and_not_pi065_n396 (not_pi065, n396, and_not_pi065_n396);
	AND2X1 g_and_pi047_n641 (n641, pi047, and_pi047_n641);
	BUFX2 g_n903 (and_pi098_pi106, n903);
	INVX1 g_not_pi003_5 (pi003, not_pi003_5);
	BUFX2 g_n1491 (and_not_n1489_not_n1490, n1491);
	INVX1 g_not_n900 (n900, not_n900);
	BUFX2 g_n371 (and_not_n368_not_n370, n371);
	BUFX2 g_po067 (po067_driver, po067);
	INVX1 g_not_n1482 (n1482, not_n1482);
	INVX1 g_not_pi138_490 (pi138, not_pi138_490);
	BUFX2 g_n390 (and_not_pi042_not_pi044, n390);
	INVX1 g_not_n1395 (n1395, not_n1395);
	INVX1 g_not_n1467 (n1467, not_n1467);
	AND2X1 g_and_not_pi129_39098210485829880490_not_n887 (not_pi129_39098210485829880490, not_n887, and_not_pi129_39098210485829880490_not_n887);
	AND2X1 g_and_n584_n650 (n584, n650, and_n584_n650);
	BUFX2 g_n983 (and_pi044_pi082, n983);
	BUFX2 g_n1484 (and_pi138_not_n1483, n1484);
	AND2X1 g_and_not_pi129_9_not_n520 (not_pi129_9, not_n520, and_not_pi129_9_not_n520);
	INVX1 g_not_n973 (n973, not_n973);
	INVX1 g_not_n875 (n875, not_n875);
	BUFX2 g_n938 (and_not_n933_n937, n938);
	INVX1 g_not_pi004_1 (pi004, not_pi004_1);
	AND2X1 g_and_not_n1064_not_n1066 (not_n1064, not_n1066, and_not_n1064_not_n1066);
	AND2X1 g_and_not_n809_not_n815 (not_n809, not_n815, and_not_n809_not_n815);
	BUFX2 g_n1508 (and_not_n1503_not_n1507, n1508);
	BUFX2 g_n849 (and_not_n846_not_n848, n849);
	AND2X1 g_and_n1049_n1054 (n1054, n1049, and_n1049_n1054);
	BUFX2 g_n907 (and_not_pi106_5_not_n906, n907);
	AND2X1 g_and_not_pi136_403536070_pi141 (pi141, not_pi136_403536070, and_not_pi136_403536070_pi141);
	INVX1 g_not_n581 (n581, not_n581);
	AND2X1 g_and_n403_n405 (n403, n405, and_n403_n405);
	BUFX2 g_n1290 (and_pi070_not_n1247_5, n1290);
	AND2X1 g_and_n856_n1223 (n1223, n856, and_n856_n1223);
	BUFX2 g_n1355 (and_not_pi137_2_not_n1354, n1355);
	BUFX2 g_n1553 (and_not_pi064_not_pi138_8235430, n1553);
	AND2X1 g_and_not_pi051_not_pi052 (not_pi052, not_pi051, and_not_pi051_not_pi052);
	INVX1 g_not_pi097_1 (pi097, not_pi097_1);
	BUFX2 g_n1438 (and_not_n1436_not_n1437, n1438);
	INVX1 g_not_pi110_3 (pi110, not_pi110_3);
	AND2X1 g_and_pi143_n1325 (n1325, pi143, and_pi143_n1325);
	INVX1 g_not_pi026_8 (pi026, not_pi026_8);
	INVX1 g_not_n1562 (n1562, not_n1562);
	INVX1 g_not_pi004_0 (pi004, not_pi004_0);
	AND2X1 g_and_n1251_n1296 (n1251, n1296, and_n1251_n1296);
	INVX1 g_not_pi008_3 (pi008, not_pi008_3);
	AND2X1 g_and_n1251_n1286 (n1251, n1286, and_n1251_n1286);
	AND2X1 g_and_pi097_not_n1423_1 (not_n1423_1, pi097, and_pi097_not_n1423_1);
	INVX1 g_not_pi027_3430 (pi027, not_pi027_3430);
	BUFX2 g_n1393 (and_not_n1391_not_n1392, n1393);
	INVX1 g_not_n1371 (n1371, not_n1371);
	BUFX2 g_n626 (and_not_pi129_8235430_not_n625, n626);
	AND2X1 g_and_not_pi005_4_n479 (n479, not_pi005_4, and_not_pi005_4_n479);
	AND2X1 g_and_not_n843_0_not_n1575 (not_n843_0, not_n1575, and_not_n843_0_not_n1575);
	BUFX2 g_n1000 (and_pi082_not_n407, n1000);
	INVX1 g_not_n1002 (n1002, not_n1002);
	BUFX2 g_po107 (po107_driver, po107);
	AND2X1 g_and_pi004_not_pi054 (not_pi054, pi004, and_pi004_not_pi054);
	INVX1 g_not_pi007_8 (pi007, not_pi007_8);
	AND2X1 g_and_not_n557_not_n564 (not_n557, not_n564, and_not_n557_not_n564);
	BUFX2 g_n1423 (and_not_n1420_not_n1422, n1423);
	INVX1 g_not_pi129_70 (pi129, not_pi129_70);
	INVX1 g_not_pi015_1 (pi015, not_pi015_1);
	AND2X1 g_and_pi008_not_pi017_3 (pi008, not_pi017_3, and_pi008_not_pi017_3);
	INVX1 g_not_pi018_3 (pi018, not_pi018_3);
	INVX1 g_not_pi027_1 (pi027, not_pi027_1);
	AND2X1 g_and_n1086_n1087 (n1087, n1086, and_n1086_n1087);
	BUFX2 g_n798 (and_not_n793_not_n797, n798);
	BUFX2 g_n328 (and_not_n325_not_n327, n328);
	BUFX2 g_n1070 (and_pi082_not_n1069, n1070);
	AND2X1 g_and_not_pi129_32199057558131797268376070_not_n961 (not_n961, not_pi129_32199057558131797268376070, and_not_pi129_32199057558131797268376070_not_n961);
	INVX1 g_not_n1320 (n1320, not_n1320);
	INVX1 g_not_pi056_0 (pi056, not_pi056_0);
	INVX1 g_not_n437 (n437, not_n437);
	AND2X1 g_and_pi021_not_pi054_24010 (not_pi054_24010, pi021, and_pi021_not_pi054_24010);
	AND2X1 g_and_pi146_n1414 (pi146, n1414, and_pi146_n1414);
	BUFX2 g_n778 (and_n762_not_n777, n778);
	INVX1 g_not_n848 (n848, not_n848);
	AND2X1 g_and_n776_n778 (n776, n778, and_n776_n778);
	BUFX2 g_n475 (and_n473_n474, n475);
	BUFX2 g_n549 (and_not_pi028_0_n548, n549);
	BUFX2 g_n763 (and_not_n728_0_n762, n763);
	AND2X1 g_and_n688_n976 (n688, n976, and_n688_n976);
	BUFX2 g_n606 (and_not_pi025_1_not_pi028_1, n606);
	BUFX2 g_po081 (po081_driver, po081);
	AND2X1 g_and_not_pi011_5_n311 (n311, not_pi011_5, and_not_pi011_5_n311);
	BUFX2 g_n698 (and_n399_n697, n698);
	BUFX2 g_n1572 (and_not_pi129_10045252112690790399992215344966975021805416861747224664747430_not_n1571, n1572);
	AND2X1 g_and_pi029_not_pi097_0 (pi029, not_pi097_0, and_pi029_not_pi097_0);
	AND2X1 g_and_not_pi129_1915812313805664144010_not_n901 (not_n901, not_pi129_1915812313805664144010, and_not_pi129_1915812313805664144010_not_n901);
	INVX1 g_not_pi116_4 (pi116, not_pi116_4);
	BUFX2 g_n767 (and_pi100_not_n766, n767);
	INVX1 g_not_n1202 (n1202, not_n1202);
	BUFX2 g_n361 (and_not_pi007_3_not_n360, n361);
	AND2X1 g_and_n369_n417 (n369, n417, and_n369_n417);
	AND2X1 g_and_n417_n598 (n417, n598, and_n417_n598);
	BUFX2 g_n1076 (and_n1073_n1075, n1076);
	BUFX2 g_n1036 (and_n385_n1035, n1036);
	BUFX2 g_po020 (po020_driver, po020);
	INVX1 g_not_n1383 (n1383, not_n1383);
	INVX1 g_not_pi027_2 (pi027, not_pi027_2);
	BUFX2 g_po061 (po061_driver, po061);
	AND2X1 g_and_not_pi116_2_not_n796 (not_n796, not_pi116_2, and_not_pi116_2_not_n796);
	AND2X1 g_and_n927_n955 (n955, n927, and_n927_n955);
	BUFX2 g_n937 (and_not_pi129_657123623635342801395430_not_n936, n937);
	BUFX2 g_n344 (and_not_pi010_0_not_pi022_0, n344);
	INVX1 g_not_pi129_3 (pi129, not_pi129_3);
	AND2X1 g_and_n568_n572 (n568, n572, and_n568_n572);
	INVX1 g_not_pi015 (pi015, not_pi015);
	AND2X1 g_and_not_n883_not_n884 (not_n884, not_n883, and_not_n883_not_n884);
	INVX1 g_not_pi136_8235430 (pi136, not_pi136_8235430);
	AND2X1 g_and_not_n1085_n1098 (not_n1085, n1098, and_not_n1085_n1098);
	INVX1 g_not_n943 (n943, not_n943);
	BUFX2 g_n1197 (and_n1192_n1196, n1197);
	BUFX2 g_n623 (and_n356_n622, n623);
	BUFX2 g_n539 (and_not_pi011_4_n418, n539);
	BUFX2 g_n1331 (and_pi143_n1325, n1331);
	BUFX2 g_po104_driver (and_not_pi129_103677930763188441902487387275962551382129494864490_not_n1393, po104_driver);
	INVX1 g_not_pi005_4 (pi005, not_pi005_4);
	INVX1 g_not_pi136 (pi136, not_pi136);
	BUFX2 g_n318 (and_not_pi013_0_not_n317, n318);
	INVX1 g_not_pi136_168070 (pi136, not_pi136_168070);
	INVX1 g_not_n983_0 (n983, not_n983_0);
	BUFX2 g_n544 (and_pi013_not_pi054_8, n544);
	AND2X1 g_and_pi141_n1325 (n1325, pi141, and_pi141_n1325);
	INVX1 g_not_n306 (n306, not_n306);
	BUFX2 g_n583 (and_not_pi045_2_n399, n583);
	BUFX2 g_po112_driver (and_not_pi129_597682638941559493067901192655856192170251494124306816490_not_n1434, po112_driver);
	INVX1 g_not_pi013_0 (pi013, not_pi013_0);
	BUFX2 g_n759 (and_not_pi129_6782230728490_not_n758, n759);
	BUFX2 g_n935 (and_pi038_n641, n935);
	AND2X1 g_and_pi100_not_n766 (not_n766, pi100, and_pi100_not_n766);
	BUFX2 g_n1262 (and_n1251_n1261, n1262);
	AND2X1 g_and_n838_n851 (n838, n851, and_n838_n851);
	BUFX2 g_n927 (and_n401_n926, n927);
	INVX1 g_not_pi129_57648010 (pi129, not_pi129_57648010);
	INVX1 g_not_n1029 (n1029, not_n1029);
	BUFX2 g_n1482 (and_pi094_n1324, n1482);
	BUFX2 g_n573 (and_n391_n572, n573);
	AND2X1 g_and_not_pi045_2_n399 (n399, not_pi045_2, and_not_pi045_2_n399);
	AND2X1 g_and_not_pi027_not_n734 (not_n734, not_pi027, and_not_pi027_not_n734);
	BUFX2 g_po041_driver (and_n772_n774, po041_driver);
	AND2X1 g_and_not_pi085_490_not_n1221 (not_pi085_490, not_n1221, and_not_pi085_490_not_n1221);
	BUFX2 g_n521 (and_not_pi129_9_not_n520, n521);
	BUFX2 g_po047 (po047_driver, po047);
	INVX1 g_not_pi021 (pi021, not_pi021);
	INVX1 g_not_pi085_3430 (pi085, not_pi085_3430);
	AND2X1 g_and_n819_n820 (n819, n820, and_n819_n820);
	BUFX2 g_n1035 (and_not_pi002_3_n399, n1035);
	BUFX2 g_po134 (po134_driver, po134);
	INVX1 g_not_n1140 (n1140, not_n1140);
	BUFX2 g_n891 (and_pi034_not_pi109_3, n891);
	BUFX2 g_n450 (and_not_pi018_0_n449, n450);
	AND2X1 g_and_not_pi026_9_not_n853 (not_pi026_9, not_n853, and_not_pi026_9_not_n853);
	INVX1 g_not_n948 (n948, not_n948);
	AND2X1 g_and_not_n1580_not_n1584 (not_n1584, not_n1580, and_not_n1580_not_n1584);
	AND2X1 g_and_n663_n666 (n663, n666, and_n663_n666);
	INVX1 g_not_pi129_4 (pi129, not_pi129_4);
	INVX1 g_not_n600 (n600, not_n600);
	AND2X1 g_and_not_pi129_152867006319425761937651857692768264010_not_n1202 (not_pi129_152867006319425761937651857692768264010, not_n1202, and_not_pi129_152867006319425761937651857692768264010_not_n1202);
	BUFX2 g_n645 (and_n640_n644, n645);
	AND2X1 g_and_not_pi085_10_n1187 (n1187, not_pi085_10, and_not_pi085_10_n1187);
	AND2X1 g_and_not_n1534_not_n1535 (not_n1535, not_n1534, and_not_n1534_not_n1535);
	AND2X1 g_and_not_pi003_0_n456 (not_pi003_0, n456, and_not_pi003_0_n456);
	BUFX2 g_n1253 (and_not_n1248_not_n1252, n1253);
	AND2X1 g_and_not_n799_n807 (not_n799, n807, and_not_n799_n807);
	AND2X1 g_and_not_n1195_not_n1197 (not_n1195, not_n1197, and_not_n1195_not_n1197);
	AND2X1 g_and_pi136_not_pi138_4 (pi136, not_pi138_4, and_pi136_not_pi138_4);
	AND2X1 g_and_pi082_not_n690 (not_n690, pi082, and_pi082_not_n690);
	INVX1 g_not_pi112 (pi112, not_pi112);
	AND2X1 g_and_not_pi137_9_not_n1542 (not_n1542, not_pi137_9, and_not_pi137_9_not_n1542);
	INVX1 g_not_n1513 (n1513, not_n1513);
	BUFX2 g_po008 (po008_driver, po008);
	AND2X1 g_and_pi085_n774 (pi085, n774, and_pi085_n774);
	BUFX2 g_n1369 (and_not_pi085_3430_not_n725_0, n1369);
	BUFX2 g_n862 (and_pi060_pi109, n862);
	AND2X1 g_and_n379_not_n966 (n379, not_n966, and_n379_not_n966);
	BUFX2 g_n531 (and_not_n523_not_n530, n531);
	BUFX2 g_po128_driver (and_not_pi003_5585458640832840070_n1598, po128_driver);
	BUFX2 g_n1167 (and_not_n1164_not_n1166, n1167);
	INVX1 g_not_n843_0 (n843, not_n843_0);
	AND2X1 g_and_pi082_not_n1089 (pi082, not_n1089, and_pi082_not_n1089);
	INVX1 g_not_pi038 (pi038, not_pi038);
	AND2X1 g_and_pi124_pi138 (pi138, pi124, and_pi124_pi138);
	INVX1 g_not_pi038_1 (pi038, not_pi038_1);
	BUFX2 g_n312 (and_not_pi007_0_pi013, n312);
	AND2X1 g_and_pi140_n1325 (n1325, pi140, and_pi140_n1325);
	INVX1 g_not_n593 (n593, not_n593);
	INVX1 g_not_n455 (n455, not_n455);
	INVX1 g_not_pi054_3430 (pi054, not_pi054_3430);
	AND2X1 g_and_not_pi129_6168735096280623662907561568153897267931784070_not_n1367 (not_pi129_6168735096280623662907561568153897267931784070, not_n1367, and_not_pi129_6168735096280623662907561568153897267931784070_not_n1367);
	INVX1 g_not_n390 (n390, not_n390);
	BUFX2 g_n1134 (and_not_n1130_n1133, n1134);
	AND2X1 g_and_not_pi129_445676403263631959001900459745680070_not_n1142 (not_pi129_445676403263631959001900459745680070, not_n1142, and_not_pi129_445676403263631959001900459745680070_not_n1142);
	AND2X1 g_and_not_pi062_not_pi138_1 (not_pi062, not_pi138_1, and_not_pi062_not_pi138_1);
	BUFX2 g_po016 (po016_driver, po016);
	INVX1 g_not_pi018 (pi018, not_pi018);
	INVX1 g_not_n595 (n595, not_n595);
	AND2X1 g_and_not_pi027_10_not_n1180 (not_pi027_10, not_n1180, and_not_pi027_10_not_n1180);
	AND2X1 g_and_n629_n632 (n629, n632, and_n629_n632);
	BUFX2 g_n479 (and_not_pi006_3_n341, n479);
	INVX1 g_not_pi029_0 (pi029, not_pi029_0);
	AND2X1 g_and_pi070_not_n1247_5 (not_n1247_5, pi070, and_pi070_not_n1247_5);
	BUFX2 g_n1349 (and_pi136_not_n1348, n1349);
	INVX1 g_not_pi129_35561530251773635572553173835655155124070416738520070 (pi129, not_pi129_35561530251773635572553173835655155124070416738520070);
	BUFX2 g_n1597 (and_not_n1594_not_n1596, n1597);
	INVX1 g_not_n565 (n565, not_n565);
	BUFX2 g_n1536 (and_not_n1534_not_n1535, n1536);
	AND2X1 g_and_n569_n570 (n569, n570, and_n569_n570);
	BUFX2 g_n517 (and_n322_n516, n517);
	INVX1 g_not_pi085_2 (pi085, not_pi085_2);
	BUFX2 g_n1057 (and_not_n379_10_not_n1056, n1057);
	AND2X1 g_and_not_n846_not_n848 (not_n848, not_n846, and_not_n846_not_n848);
	INVX1 g_not_pi012_4 (pi012, not_pi012_4);
	BUFX2 g_n1250 (and_not_pi140_n1249, n1250);
	AND2X1 g_and_not_pi129_225393402906922580878632490_not_n979 (not_n979, not_pi129_225393402906922580878632490, and_not_pi129_225393402906922580878632490_not_n979);
	AND2X1 g_and_pi078_not_n1325 (not_n1325, pi078, and_pi078_not_n1325);
	INVX1 g_not_pi116 (pi116, not_pi116);
	BUFX2 g_n1023 (and_not_n1019_not_n1022, n1023);
	AND2X1 g_and_pi032_pi136 (pi136, pi032, and_pi032_pi136);
	AND2X1 g_and_not_pi003_6782230728490_n1210 (n1210, not_pi003_6782230728490, and_not_pi003_6782230728490_n1210);
	BUFX2 g_n314 (and_not_pi007_1_n311, n314);
	AND2X1 g_and_not_n1164_0_not_n1170 (not_n1170, not_n1164_0, and_not_n1164_0_not_n1170);
	AND2X1 g_and_pi002_not_n412 (pi002, not_n412, and_pi002_not_n412);
	BUFX2 g_n915 (and_not_n910_not_n914, n915);
	INVX1 g_not_n782 (n782, not_n782);
	INVX1 g_not_pi043_3 (pi043, not_pi043_3);
	AND2X1 g_and_n487_n667 (n487, n667, and_n487_n667);
	BUFX2 g_n322 (and_not_pi013_1_pi014, n322);
	INVX1 g_not_pi136_0 (pi136, not_pi136_0);
	INVX1 g_not_n1138 (n1138, not_n1138);
	BUFX2 g_po112 (po112_driver, po112);
	BUFX2 g_n1276 (and_pi067_not_n1271_0, n1276);
	INVX1 g_not_pi129_968890104070 (pi129, not_pi129_968890104070);
	AND2X1 g_and_not_pi003_113988951853731430_n1572 (n1572, not_pi003_113988951853731430, and_not_pi003_113988951853731430_n1572);
	INVX1 g_not_pi049 (pi049, not_pi049);
	INVX1 g_not_pi138_9 (pi138, not_pi138_9);
	BUFX2 g_n764 (and_not_pi096_0_n763, n764);
	AND2X1 g_and_not_n321_not_n323 (not_n323, not_n321, and_not_n321_not_n323);
	AND2X1 g_and_not_pi115_pi138 (not_pi115, pi138, and_not_pi115_pi138);
	AND2X1 g_and_not_n1359_not_n1361 (not_n1361, not_n1359, and_not_n1359_not_n1361);
	INVX1 g_not_pi013_4 (pi013, not_pi013_4);
	INVX1 g_not_n379_0 (n379, not_n379_0);
	INVX1 g_not_pi005_2 (pi005, not_pi005_2);
	INVX1 g_not_n313 (n313, not_n313);
	BUFX2 g_po102 (po102_driver, po102);
	AND2X1 g_and_not_pi129_7_not_n495 (not_n495, not_pi129_7, and_not_pi129_7_not_n495);
	AND2X1 g_and_pi067_not_n379_8 (pi067, not_n379_8, and_pi067_not_n379_8);
	BUFX2 g_n440 (and_pi005_not_pi054_0, n440);
	BUFX2 g_n445 (and_not_pi013_4_n417, n445);
	AND2X1 g_and_pi097_pi116 (pi116, pi097, and_pi097_pi116);
	BUFX2 g_n743 (and_not_pi026_0_not_pi085_1, n743);
	INVX1 g_not_n669 (n669, not_n669);
	INVX1 g_not_pi129_7 (pi129, not_pi129_7);
	AND2X1 g_and_not_pi146_0_n1271 (n1271, not_pi146_0, and_not_pi146_0_n1271);
	AND2X1 g_and_not_pi137_70_pi138 (pi138, not_pi137_70, and_not_pi137_70_pi138);
	INVX1 g_not_n886 (n886, not_n886);
	AND2X1 g_and_not_pi106_6_not_n913 (not_pi106_6, not_n913, and_not_pi106_6_not_n913);
	AND2X1 g_and_not_n1436_not_n1437 (not_n1436, not_n1437, and_not_n1436_not_n1437);
	BUFX2 g_n395 (and_pi082_not_n394, n395);
	INVX1 g_not_n362 (n362, not_n362);
	BUFX2 g_n1026 (and_n399_n704, n1026);
	INVX1 g_not_pi140 (pi140, not_pi140);
	INVX1 g_not_n1027 (n1027, not_n1027);
	BUFX2 g_n1018 (and_n927_n1017, n1018);
	BUFX2 g_n1085 (and_not_pi048_3_not_n1084, n1085);
	AND2X1 g_and_not_n1072_n1077 (not_n1072, n1077, and_not_n1072_n1077);
	BUFX2 g_n1168 (and_pi094_not_n1167, n1168);
	INVX1 g_not_n738_0 (n738, not_n738_0);
	AND2X1 g_and_pi058_not_pi116_7 (not_pi116_7, pi058, and_pi058_not_pi116_7);
	INVX1 g_not_n1176 (n1176, not_n1176);
	AND2X1 g_and_not_pi003_8235430_n771 (n771, not_pi003_8235430, and_not_pi003_8235430_n771);
	AND2X1 g_and_pi031_n1360 (n1360, pi031, and_pi031_n1360);
	AND2X1 g_and_pi084_not_n1325_4 (pi084, not_n1325_4, and_pi084_not_n1325_4);
	INVX1 g_not_n1403 (n1403, not_n1403);
	BUFX2 g_po079_driver (or_pi129_n1263, po079_driver);
	BUFX2 g_n1172 (and_not_n1169_not_n1171, n1172);
	INVX1 g_not_n427 (n427, not_n427);
	INVX1 g_not_pi110_4 (pi110, not_pi110_4);
	AND2X1 g_and_n291_n676 (n676, n291, and_n291_n676);
	AND2X1 g_and_pi029_pi110 (pi029, pi110, and_pi029_pi110);
	INVX1 g_not_pi019_1 (pi019, not_pi019_1);
	INVX1 g_not_pi003_47475615099430 (pi003, not_pi003_47475615099430);
	AND2X1 g_and_pi025_not_n726 (not_n726, pi025, and_pi025_not_n726);
	BUFX2 g_n1224 (and_pi085_n787, n1224);
	INVX1 g_not_n1332 (n1332, not_n1332);
	BUFX2 g_po070_driver (and_not_po129_n1162, po070_driver);
	BUFX2 g_n741 (and_n723_n727, n741);
	BUFX2 g_n797 (and_not_pi116_2_not_n796, n797);
	BUFX2 g_n1019 (and_pi082_not_n1018, n1019);
	BUFX2 g_po061_driver (and_not_n1053_n1062, po061_driver);
	INVX1 g_not_n1501 (n1501, not_n1501);
	BUFX2 g_n635 (and_not_n628_not_n634, n635);
	INVX1 g_not_n601 (n601, not_n601);
	INVX1 g_not_n436 (n436, not_n436);
	INVX1 g_not_pi012_3 (pi012, not_pi012_3);
	INVX1 g_not_n933 (n933, not_n933);
	AND2X1 g_and_n389_n948 (n389, n948, and_n389_n948);
	INVX1 g_not_pi129_77309937197074445241370944070 (pi129, not_pi129_77309937197074445241370944070);
	AND2X1 g_and_pi082_not_n408 (not_n408, pi082, and_pi082_not_n408);
	AND2X1 g_and_not_pi129_367033682172941254412302110320336601888010_not_n1328 (not_pi129_367033682172941254412302110320336601888010, not_n1328, and_not_pi129_367033682172941254412302110320336601888010_not_n1328);
	INVX1 g_not_pi129_10 (pi129, not_pi129_10);
	BUFX2 g_n756 (and_n754_n755, n756);
	INVX1 g_not_pi129_3430 (pi129, not_pi129_3430);
	AND2X1 g_and_pi031_not_pi109_0 (not_pi109_0, pi031, and_pi031_not_pi109_0);
	INVX1 g_not_n876 (n876, not_n876);
	INVX1 g_not_n1018 (n1018, not_n1018);
	BUFX2 g_n1120 (and_n704_n1035, n1120);
	INVX1 g_not_n1595 (n1595, not_n1595);
	BUFX2 g_po074 (po074_driver, po074);
	INVX1 g_not_n411 (n411, not_n411);
	INVX1 g_not_n1247_4 (n1247, not_n1247_4);
	INVX1 g_not_pi137_10 (pi137, not_pi137_10);
	INVX1 g_not_pi145_0 (pi145, not_pi145_0);
	INVX1 g_not_pi136_490 (pi136, not_pi136_490);
	BUFX2 g_n1433 (and_pi145_n1414, n1433);
	AND2X1 g_and_pi082_not_n1001 (not_n1001, pi082, and_pi082_not_n1001);
	BUFX2 g_n1537 (and_pi136_not_n1536, n1537);
	AND2X1 g_and_n399_n697 (n399, n697, and_n399_n697);
	BUFX2 g_n577 (and_not_n379_0_not_n576, n577);
	BUFX2 g_n758 (and_not_n753_not_n757, n758);
	INVX1 g_not_n1328 (n1328, not_n1328);
	AND2X1 g_and_n819_n824 (n819, n824, and_n819_n824);
	BUFX2 g_po090 (po090_driver, po090);
	AND2X1 g_and_n311_n312 (n311, n312, and_n311_n312);
	INVX1 g_not_n1037 (n1037, not_n1037);
	INVX1 g_not_pi071 (pi071, not_pi071);
	INVX1 g_not_pi129_2824752490 (pi129, not_pi129_2824752490);
	BUFX2 g_n1056 (and_pi082_not_n1055, n1056);
	INVX1 g_not_pi054_70 (pi054, not_pi054_70);
	INVX1 g_not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430 (pi129, not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430);
	AND2X1 g_and_not_n1010_n1014 (not_n1010, n1014, and_not_n1010_n1014);
	BUFX2 g_po018_driver (and_not_pi129_2_not_n428, po018_driver);
	OR2X1 g_or_pi129_n1253 (pi129, n1253, or_pi129_n1253);
	BUFX2 g_n1271 (and_n1251_n1270, n1271);
	AND2X1 g_and_not_n365_not_n366 (not_n365, not_n366, and_not_n365_not_n366);
	BUFX2 g_n1571 (and_not_n794_0_not_n1570, n1571);
	BUFX2 g_n1194 (and_not_n1191_not_n1193, n1194);
	INVX1 g_not_n1081 (n1081, not_n1081);
	INVX1 g_not_n1338 (n1338, not_n1338);
	BUFX2 g_n538 (and_n536_n537, n538);
	AND2X1 g_and_n736_n940 (n940, n736, and_n736_n940);
	BUFX2 g_n998 (and_not_n995_n997, n998);
	INVX1 g_not_n1511 (n1511, not_n1511);
	INVX1 g_not_n917 (n917, not_n917);
	BUFX2 g_n570 (and_not_pi045_1_n384, n570);
	OR2X1 g_or_pi129_n1278 (pi129, n1278, or_pi129_n1278);
	INVX1 g_not_pi129_9 (pi129, not_pi129_9);
	INVX1 g_not_n423 (n423, not_n423);
	INVX1 g_not_pi050_2 (pi050, not_pi050_2);
	INVX1 g_not_n1386_6 (n1386, not_n1386_6);
	AND2X1 g_and_n448_n476 (n476, n448, and_n448_n476);
	INVX1 g_not_n1487 (n1487, not_n1487);
	AND2X1 g_and_not_pi003_2824752490_n859 (not_pi003_2824752490, n859, and_not_pi003_2824752490_n859);
	AND2X1 g_and_n391_n572 (n391, n572, and_n391_n572);
	AND2X1 g_and_pi061_n686 (pi061, n686, and_pi061_n686);
	BUFX2 g_n1180 (and_not_n1178_not_n1179, n1180);
	INVX1 g_not_pi003_16284135979104490 (pi003, not_pi003_16284135979104490);
	BUFX2 g_n1248 (and_pi062_not_n1247, n1248);
	BUFX2 g_n1615 (and_n549_n1614, n1615);
	AND2X1 g_and_not_pi129_4183778472590916451475308348590993345191760458870147715430_not_n1438 (not_pi129_4183778472590916451475308348590993345191760458870147715430, not_n1438, and_not_pi129_4183778472590916451475308348590993345191760458870147715430_not_n1438);
	INVX1 g_not_n715 (n715, not_n715);
	AND2X1 g_and_not_n983_not_n987 (not_n987, not_n983, and_not_n983_not_n987);
	BUFX2 g_n1544 (and_pi036_n1360, n1544);
	AND2X1 g_and_not_pi136_3430_not_n1523 (not_n1523, not_pi136_3430, and_not_pi136_3430_not_n1523);
	AND2X1 g_and_not_n730_not_n731 (not_n731, not_n730, and_not_n730_not_n731);
	BUFX2 g_n493 (and_n490_n492, n493);
	INVX1 g_not_pi003_968890104070 (pi003, not_pi003_968890104070);
	INVX1 g_not_pi003_168070 (pi003, not_pi003_168070);
	AND2X1 g_and_n642_n643 (n643, n642, and_n642_n643);
	BUFX2 g_n1356 (and_not_pi115_pi138, n1356);
	BUFX2 g_po065 (po065_driver, po065);
	INVX1 g_not_n494 (n494, not_n494);
	BUFX2 g_n1334 (and_pi080_not_n1325_1, n1334);
	AND2X1 g_and_not_pi013_3_not_n364 (not_pi013_3, not_n364, and_not_pi013_3_not_n364);
	INVX1 g_not_n495 (n495, not_n495);
	AND2X1 g_and_not_pi136_490_not_n1517 (not_n1517, not_pi136_490, and_not_pi136_490_not_n1517);
	BUFX2 g_po021_driver (and_not_pi003_1_n470, po021_driver);
	AND2X1 g_and_not_n1538_not_n1539 (not_n1539, not_n1538, and_not_n1538_not_n1539);
	INVX1 g_not_n852 (n852, not_n852);
	INVX1 g_not_n1389 (n1389, not_n1389);
	INVX1 g_not_pi045 (pi045, not_pi045);
	AND2X1 g_and_not_n534_not_n540 (not_n534, not_n540, and_not_n534_not_n540);
	AND2X1 g_and_pi136_not_n1348 (not_n1348, pi136, and_pi136_not_n1348);
	INVX1 g_not_n1498 (n1498, not_n1498);
	BUFX2 g_n1078 (and_not_n1072_n1077, n1078);
	INVX1 g_not_n335 (n335, not_n335);
	BUFX2 g_n1292 (and_n1251_n1291, n1292);
	INVX1 g_not_pi026_7 (pi026, not_pi026_7);
	AND2X1 g_and_not_pi112_n1324 (not_pi112, n1324, and_not_pi112_n1324);
	INVX1 g_not_n648 (n648, not_n648);
	AND2X1 g_and_not_n1058_n1061 (n1061, not_n1058, and_not_n1058_n1061);
	INVX1 g_not_n1230 (n1230, not_n1230);
	AND2X1 g_and_not_n379_4_not_n957 (not_n379_4, not_n957, and_not_n379_4_not_n957);
	AND2X1 g_and_not_pi129_138412872010_not_n685 (not_n685, not_pi129_138412872010, and_not_pi129_138412872010_not_n685);
	INVX1 g_not_pi048_3 (pi048, not_pi048_3);
	BUFX2 g_n562 (and_n344_n561, n562);
	BUFX2 g_n847 (and_pi027_n838, n847);
	BUFX2 g_n639 (and_not_pi024_1_n380, n639);
	BUFX2 g_n1523 (and_not_n1521_not_n1522, n1523);
	INVX1 g_not_pi021_2 (pi021, not_pi021_2);
	BUFX2 g_po063_driver (and_not_n1085_n1098, po063_driver);
	INVX1 g_not_pi003_403536070 (pi003, not_pi003_403536070);
	AND2X1 g_and_pi137_not_n1526 (pi137, not_n1526, and_pi137_not_n1526);
	INVX1 g_not_pi051 (pi051, not_pi051);
	INVX1 g_not_n988 (n988, not_n988);
	INVX1 g_not_n544 (n544, not_n544);
	AND2X1 g_and_not_pi009_5_not_pi010_3 (not_pi009_5, not_pi010_3, and_not_pi009_5_not_pi010_3);
	AND2X1 g_and_not_pi129_103677930763188441902487387275962551382129494864490_not_n1393 (not_pi129_103677930763188441902487387275962551382129494864490, not_n1393, and_not_pi129_103677930763188441902487387275962551382129494864490_not_n1393);
	AND2X1 g_and_not_n1342_not_n1343 (not_n1342, not_n1343, and_not_n1342_not_n1343);
	BUFX2 g_po023 (po023_driver, po023);
	AND2X1 g_and_pi082_n1582 (n1582, pi082, and_pi082_n1582);
	BUFX2 g_n1281 (and_not_pi141_n1249, n1281);
	AND2X1 g_and_n448_n631 (n631, n448, and_n448_n631);
	AND2X1 g_and_not_pi116_9_n1192 (not_pi116_9, n1192, and_not_pi116_9_n1192);
	BUFX2 g_n1330 (and_pi079_not_n1325_0, n1330);
	INVX1 g_not_n883 (n883, not_n883);
	BUFX2 g_n501 (and_n332_n500, n501);
	AND2X1 g_and_not_n975_n980 (not_n975, n980, and_not_n975_n980);
	BUFX2 g_n911 (and_pi036_pi109, n911);
	BUFX2 g_n578 (and_not_pi070_n577, n578);
	BUFX2 g_n676 (and_not_pi009_5_not_pi010_3, n676);
	AND2X1 g_and_not_pi129_10045252112690790399992215344966975021805416861747224664747430_not_n1571 (not_n1571, not_pi129_10045252112690790399992215344966975021805416861747224664747430, and_not_pi129_10045252112690790399992215344966975021805416861747224664747430_not_n1571);
	INVX1 g_not_n809 (n809, not_n809);
	BUFX2 g_n1547 (and_not_n1545_not_n1546, n1547);
	AND2X1 g_and_pi022_not_pi054_168070 (not_pi054_168070, pi022, and_pi022_not_pi054_168070);
	AND2X1 g_and_not_n1019_not_n1022 (not_n1022, not_n1019, and_not_n1019_not_n1022);
	BUFX2 g_po011_driver (pi000, po011_driver);
	AND2X1 g_and_n390_n403 (n403, n390, and_n390_n403);
	INVX1 g_not_n1346 (n1346, not_n1346);
	AND2X1 g_and_not_pi043_2_n387 (not_pi043_2, n387, and_not_pi043_2_n387);
	INVX1 g_not_pi053_1 (pi053, not_pi053_1);
	INVX1 g_not_n540 (n540, not_n540);
	INVX1 g_not_pi138_6 (pi138, not_pi138_6);
	BUFX2 g_n1372 (and_not_n761_0_not_n1371, n1372);
	INVX1 g_not_n766 (n766, not_n766);
	INVX1 g_not_pi021_3 (pi021, not_pi021_3);
	BUFX2 g_po111 (po111_driver, po111);
	AND2X1 g_and_not_pi129_273687473400809163430_not_n894 (not_pi129_273687473400809163430, not_n894, and_not_pi129_273687473400809163430_not_n894);
	AND2X1 g_and_not_pi027_490_not_n1226 (not_n1226, not_pi027_490, and_not_pi027_490_not_n1226);
	INVX1 g_not_pi054_8235430 (pi054, not_pi054_8235430);
	BUFX2 g_po010_driver (pi001, po010_driver);
	BUFX2 g_n1324 (and_not_pi136_0_pi137, n1324);
	INVX1 g_not_n1512 (n1512, not_n1512);
	INVX1 g_not_n804 (n804, not_n804);
	AND2X1 g_and_pi064_n1071 (pi064, n1071, and_pi064_n1071);
	INVX1 g_not_pi129_1915812313805664144010 (pi129, not_pi129_1915812313805664144010);
	INVX1 g_not_pi026_2 (pi026, not_pi026_2);
	INVX1 g_not_n863 (n863, not_n863);
	BUFX2 g_n655 (and_pi002_n645, n655);
	AND2X1 g_and_not_pi039_n722 (n722, not_pi039, and_not_pi039_n722);
	INVX1 g_not_n718 (n718, not_n718);
	AND2X1 g_and_pi028_not_n798 (pi028, not_n798, and_pi028_not_n798);
	AND2X1 g_and_pi028_n442 (pi028, n442, and_pi028_n442);
	BUFX2 g_n979 (and_n976_n978, n979);
	AND2X1 g_and_not_pi015_0_n573 (n573, not_pi015_0, and_not_pi015_0_n573);
	BUFX2 g_n786 (and_not_pi003_57648010_n785, n786);
	OR2X1 g_or_pi129_n1159 (pi129, n1159, or_pi129_n1159);
	BUFX2 g_n1265 (and_pi065_not_n1247_2, n1265);
	BUFX2 g_n1594 (and_not_pi054_1176490_not_pi113_0, n1594);
	BUFX2 g_n350 (and_n343_n349, n350);
	AND2X1 g_and_not_pi027_1_not_pi085_3 (not_pi027_1, not_pi085_3, and_not_pi027_1_not_pi085_3);
	BUFX2 g_n1147 (and_n724_n1146, n1147);
	AND2X1 g_and_n1192_n1200 (n1192, n1200, and_n1192_n1200);
	INVX1 g_not_n1080 (n1080, not_n1080);
	AND2X1 g_and_n301_not_n328 (not_n328, n301, and_n301_not_n328);
	AND2X1 g_and_n724_n1146 (n724, n1146, and_n724_n1146);
	AND2X1 g_and_not_pi027_3_n713 (n713, not_pi027_3, and_not_pi027_3_n713);
	INVX1 g_not_n921 (n921, not_n921);
	BUFX2 g_n1606 (and_not_pi004_2_not_pi012_6, n1606);
	AND2X1 g_and_not_n718_not_n738 (not_n718, not_n738, and_not_n718_not_n738);
	INVX1 g_not_n1423_1 (n1423, not_n1423_1);
	AND2X1 g_and_not_pi129_70_not_n541 (not_n541, not_pi129_70, and_not_pi129_70_not_n541);
	INVX1 g_not_n1352 (n1352, not_n1352);
	INVX1 g_not_n910 (n910, not_n910);
	BUFX2 g_po107_driver (and_not_pi129_35561530251773635572553173835655155124070416738520070_not_n1405, po107_driver);
	AND2X1 g_and_not_pi003_6_n532 (n532, not_pi003_6, and_not_pi003_6_n532);
	BUFX2 g_n766 (and_not_n764_not_n765, n766);
	BUFX2 g_n1450 (and_not_n1448_not_n1449, n1450);
	AND2X1 g_and_not_pi139_n1249 (not_pi139, n1249, and_not_pi139_n1249);
	BUFX2 g_n1515 (and_pi125_pi138, n1515);
	BUFX2 g_n859 (and_not_pi129_16284135979104490_not_n858, n859);
	INVX1 g_not_n507 (n507, not_n507);
	INVX1 g_not_n1287 (n1287, not_n1287);
	AND2X1 g_and_pi036_n1360 (pi036, n1360, and_pi036_n1360);
	AND2X1 g_and_not_pi129_1742514982336908143055105517947102601079450420187483430_not_n1417 (not_n1417, not_pi129_1742514982336908143055105517947102601079450420187483430, and_not_pi129_1742514982336908143055105517947102601079450420187483430_not_n1417);
	INVX1 g_not_n1539 (n1539, not_n1539);
	BUFX2 g_po045_driver (and_not_pi129_113988951853731430_not_n866, po045_driver);
	AND2X1 g_and_n927_n1006 (n1006, n927, and_n927_n1006);
	BUFX2 g_n305 (and_n297_n304, n305);
	BUFX2 g_n1437 (and_pi145_n1386, n1437);
	BUFX2 g_n1175 (and_not_pi026_490_pi037, n1175);
	AND2X1 g_and_not_n1205_not_n1208 (not_n1208, not_n1205, and_not_n1205_not_n1208);
	AND2X1 g_and_n379_not_n986 (n379, not_n986, and_n379_not_n986);
	INVX1 g_not_n1546 (n1546, not_n1546);
	INVX1 g_not_pi026_6 (pi026, not_pi026_6);
	BUFX2 g_n1610 (and_not_pi003_39098210485829880490_n1609, n1610);
	BUFX2 g_n1595 (and_not_pi011_6_not_pi022_4, n1595);
	INVX1 g_not_pi053_0 (pi053, not_pi053_0);
	BUFX2 g_n1489 (and_not_pi063_pi136, n1489);
	AND2X1 g_and_pi085_pi116 (pi085, pi116, and_pi085_pi116);
	INVX1 g_not_pi026_3430 (pi026, not_pi026_3430);
	AND2X1 g_and_pi080_not_pi138_3430 (not_pi138_3430, pi080, and_pi080_not_pi138_3430);
	BUFX2 g_n1500 (and_not_pi068_pi136, n1500);
	AND2X1 g_and_not_pi129_not_n338 (not_n338, not_pi129, and_not_pi129_not_n338);
	BUFX2 g_n990 (and_not_pi044_2_n649, n990);
	BUFX2 g_n1616 (and_not_n1613_not_n1615, n1616);
	BUFX2 g_po098_driver (or_n1355_n1363, po098_driver);
	INVX1 g_not_pi142_0 (pi142, not_pi142_0);
	BUFX2 g_n346 (and_not_pi005_0_not_pi006_1, n346);
	INVX1 g_not_pi129_1070069044235980333563563003849377848070 (pi129, not_pi129_1070069044235980333563563003849377848070);
	BUFX2 g_n1415 (and_pi094_not_n1414, n1415);
	AND2X1 g_and_not_pi012_n295 (not_pi012, n295, and_not_pi012_n295);
	BUFX2 g_n845 (and_not_n842_not_n844, n845);
	BUFX2 g_n836 (and_not_pi058_3_not_n835, n836);
	AND2X1 g_and_n379_not_n950 (not_n950, n379, and_n379_not_n950);
	BUFX2 g_n974 (and_not_n379_5_not_n973, n974);
	AND2X1 g_and_not_pi005_2_n450 (n450, not_pi005_2, and_not_pi005_2_n450);
	BUFX2 g_n680 (and_n677_n679, n680);
	BUFX2 g_n1375 (and_n774_n1374, n1375);
	AND2X1 g_and_not_n1594_not_n1596 (not_n1594, not_n1596, and_not_n1594_not_n1596);
	INVX1 g_not_n1049 (n1049, not_n1049);
	AND2X1 g_and_n934_n1042 (n934, n1042, and_n934_n1042);
	AND2X1 g_and_n356_n622 (n622, n356, and_n356_n622);
	AND2X1 g_and_not_pi129_405362155971443868320658661090166738008752222510120837461924544480010_not_n1620 (not_n1620, not_pi129_405362155971443868320658661090166738008752222510120837461924544480010, and_not_pi129_405362155971443868320658661090166738008752222510120837461924544480010_not_n1620);
	BUFX2 g_n667 (and_n663_n666, n667);
	BUFX2 g_n1029 (and_pi082_not_n1028, n1029);
	INVX1 g_not_pi027_490 (pi027, not_pi027_490);
	BUFX2 g_n1555 (and_pi136_not_n1554, n1555);
	AND2X1 g_and_not_pi129_6782230728490_not_n758 (not_n758, not_pi129_6782230728490, and_not_pi129_6782230728490_not_n758);
	BUFX2 g_n1446 (and_not_n1444_not_n1445, n1446);
	AND2X1 g_and_not_pi003_5585458640832840070_n1598 (not_pi003_5585458640832840070, n1598, and_not_pi003_5585458640832840070_n1598);
	AND2X1 g_and_n990_n1105 (n1105, n990, and_n990_n1105);
	INVX1 g_not_n850 (n850, not_n850);
	AND2X1 g_and_not_n1474_not_n1475 (not_n1475, not_n1474, and_not_n1474_not_n1475);
	BUFX2 g_n1440 (and_pi099_not_n1386_6, n1440);
	INVX1 g_not_pi138_168070 (pi138, not_pi138_168070);
	BUFX2 g_n359 (and_not_n357_not_n358, n359);
	AND2X1 g_and_not_pi007_3_not_n360 (not_pi007_3, not_n360, and_not_pi007_3_not_n360);
	AND2X1 g_and_pi137_not_n1472 (pi137, not_n1472, and_pi137_not_n1472);
	AND2X1 g_and_n503_n505 (n503, n505, and_n503_n505);
	INVX1 g_not_pi013 (pi013, not_pi013);
	INVX1 g_not_n1444 (n1444, not_n1444);
	AND2X1 g_and_not_n379_0_not_n576 (not_n576, not_n379_0, and_not_n379_0_not_n576);
	AND2X1 g_and_not_pi017_4_not_pi018_2 (not_pi017_4, not_pi018_2, and_not_pi017_4_not_pi018_2);
	INVX1 g_not_pi050_4 (pi050, not_pi050_4);
	BUFX2 g_po083 (po083_driver, po083);
	INVX1 g_not_n791 (n791, not_n791);
	INVX1 g_not_n534 (n534, not_n534);
	INVX1 g_not_n1507 (n1507, not_n1507);
	BUFX2 g_n1123 (and_n379_not_n1122, n1123);
	BUFX2 g_n1050 (and_pi082_not_n1049, n1050);
	INVX1 g_not_n1008 (n1008, not_n1008);
	BUFX2 g_n1462 (and_not_pi136_5_not_n1461, n1462);
	AND2X1 g_and_pi072_n994 (pi072, n994, and_pi072_n994);
	BUFX2 g_po043_driver (and_not_pi003_403536070_n827, po043_driver);
	BUFX2 g_n1332 (and_not_n1330_not_n1331, n1332);
	AND2X1 g_and_not_pi007_7_n417 (not_pi007_7, n417, and_not_pi007_7_n417);
	AND2X1 g_and_n1073_n1075 (n1073, n1075, and_n1073_n1075);
	INVX1 g_not_n1367 (n1367, not_n1367);
	OR2X1 g_or_pi129_n1298 (pi129, n1298, or_pi129_n1298);
	AND2X1 g_and_not_pi129_2569235775210588780886114772242356213216070_not_n1332 (not_n1332, not_pi129_2569235775210588780886114772242356213216070, and_not_pi129_2569235775210588780886114772242356213216070_not_n1332);
	AND2X1 g_and_n464_n467 (n464, n467, and_n464_n467);
	INVX1 g_not_n523 (n523, not_n523);
	INVX1 g_not_n1272 (n1272, not_n1272);
	AND2X1 g_and_n515_n562 (n562, n515, and_n515_n562);
	BUFX2 g_n975 (and_pi076_n974, n975);
	INVX1 g_not_pi129_2569235775210588780886114772242356213216070 (pi129, not_pi129_2569235775210588780886114772242356213216070);
	INVX1 g_not_n321 (n321, not_n321);
	INVX1 g_not_n1372 (n1372, not_n1372);
	BUFX2 g_po110 (po110_driver, po110);
	AND2X1 g_and_not_pi110_5_n1369 (n1369, not_pi110_5, and_not_pi110_5_n1369);
	BUFX2 g_n751 (and_n748_n750, n751);
	BUFX2 g_n689 (and_n380_n688, n689);
	BUFX2 g_n1058 (and_pi075_n1057, n1058);
	INVX1 g_not_n1461 (n1461, not_n1461);
	AND2X1 g_and_not_pi129_70316764788835532799945507414768825152637918032230572653232010_not_n1576 (not_n1576, not_pi129_70316764788835532799945507414768825152637918032230572653232010, and_not_pi129_70316764788835532799945507414768825152637918032230572653232010_not_n1576);
	BUFX2 g_po033 (po033_driver, po033);
	INVX1 g_not_pi129 (pi129, not_pi129);
	BUFX2 g_n1231 (and_not_pi026_24010_not_n1230, n1231);
	BUFX2 g_po030 (po030_driver, po030);
	AND2X1 g_and_not_pi063_pi136 (not_pi063, pi136, and_not_pi063_pi136);
	BUFX2 g_n372 (and_n300_not_n371, n372);
	INVX1 g_not_n557 (n557, not_n557);
	BUFX2 g_po099_driver (and_not_pi129_6168735096280623662907561568153897267931784070_not_n1367, po099_driver);
	AND2X1 g_and_n1250_n1251 (n1251, n1250, and_n1250_n1251);
	INVX1 g_not_n815 (n815, not_n815);
	BUFX2 g_n1302 (and_not_n1300_not_n1301, n1302);
	INVX1 g_not_n1316 (n1316, not_n1316);
	BUFX2 g_n861 (and_pi030_not_pi109, n861);
	BUFX2 g_n455 (and_not_n440_not_n454, n455);
	BUFX2 g_n723 (and_not_pi039_n722, n723);
	BUFX2 g_n894 (and_not_n889_not_n893, n894);
	AND2X1 g_and_pi136_pi137 (pi137, pi136, and_pi136_pi137);
	AND2X1 g_and_not_n890_not_n891 (not_n890, not_n891, and_not_n890_not_n891);
	INVX1 g_not_n794 (n794, not_n794);
	AND2X1 g_and_n638_n990 (n638, n990, and_n638_n990);
	AND2X1 g_and_not_n1222_not_n1225 (not_n1225, not_n1222, and_not_n1222_not_n1225);
	AND2X1 g_and_not_pi096_0_n763 (not_pi096_0, n763, and_not_pi096_0_n763);
	BUFX2 g_n735 (and_not_pi027_not_n734, n735);
	AND2X1 g_and_not_pi129_5_not_n469 (not_n469, not_pi129_5, and_not_pi129_5_not_n469);
	BUFX2 g_n1475 (and_not_pi066_not_pi136_7, n1475);
	AND2X1 g_and_not_pi003_24010_n670 (n670, not_pi003_24010, and_not_pi003_24010_n670);
	AND2X1 g_and_not_n379_3430_not_n1102 (not_n1102, not_n379_3430, and_not_n379_3430_not_n1102);
	BUFX2 g_n1400 (and_pi143_n1386, n1400);
	BUFX2 g_n770 (and_not_n767_not_n769, n770);
	INVX1 g_not_pi003_4 (pi003, not_pi003_4);
	INVX1 g_not_n1508 (n1508, not_n1508);
	INVX1 g_not_pi059 (pi059, not_pi059);
	BUFX2 g_n364 (and_not_n362_not_n363, n364);
	AND2X1 g_and_n488_n489 (n489, n488, and_n488_n489);
	BUFX2 g_po004_driver (pi102, po004_driver);
	BUFX2 g_n788 (and_not_pi026_3_n787, n788);
	AND2X1 g_and_not_pi129_403536070_not_n660 (not_pi129_403536070, not_n660, and_not_pi129_403536070_not_n660);
	INVX1 g_not_n486 (n486, not_n486);
	INVX1 g_not_n425 (n425, not_n425);
	OR2X1 g_or_pi129_n1263 (n1263, pi129, or_pi129_n1263);
	INVX1 g_not_n729 (n729, not_n729);
	BUFX2 g_n1576 (and_not_n843_0_not_n1575, n1576);
	INVX1 g_not_n1348 (n1348, not_n1348);
	INVX1 g_not_n949 (n949, not_n949);
	BUFX2 g_n682 (and_not_n672_not_n681, n682);
	INVX1 g_not_pi017_3 (pi017, not_pi017_3);
	INVX1 g_not_n1517 (n1517, not_n1517);
	AND2X1 g_and_not_n755_not_n843 (not_n843, not_n755, and_not_n755_not_n843);
	AND2X1 g_and_not_pi008_2_not_pi017_2 (not_pi008_2, not_pi017_2, and_not_pi008_2_not_pi017_2);
	AND2X1 g_and_not_pi053_6_not_n1173 (not_n1173, not_pi053_6, and_not_pi053_6_not_n1173);
	AND2X1 g_and_n503_n559 (n559, n503, and_n503_n559);
	AND2X1 g_and_not_pi129_113988951853731430_not_n866 (not_n866, not_pi129_113988951853731430, and_not_pi129_113988951853731430_not_n866);
	INVX1 g_not_n1488 (n1488, not_n1488);
	AND2X1 g_and_not_pi077_not_pi138_5 (not_pi077, not_pi138_5, and_not_pi077_not_pi138_5);
	AND2X1 g_and_not_pi011_6_not_pi022_4 (not_pi022_4, not_pi011_6, and_not_pi011_6_not_pi022_4);
	AND2X1 g_and_not_pi129_4599865365447399609768010_not_n945 (not_pi129_4599865365447399609768010, not_n945, and_not_pi129_4599865365447399609768010_not_n945);
	BUFX2 g_n1293 (and_not_n1290_not_n1292, n1293);
	BUFX2 g_n491 (and_not_pi008_3_n449, n491);
	BUFX2 g_n1556 (and_pi120_pi138, n1556);
	BUFX2 g_n356 (and_n294_n355, n356);
	AND2X1 g_and_not_n713_0_not_n1530 (not_n713_0, not_n1530, and_not_n713_0_not_n1530);
	INVX1 g_not_n1082 (n1082, not_n1082);
	BUFX2 g_n818 (and_not_pi027_8_pi028, n818);
	AND2X1 g_and_not_pi065_0_not_pi138_6 (not_pi065_0, not_pi138_6, and_not_pi065_0_not_pi138_6);
	INVX1 g_not_n1407 (n1407, not_n1407);
	BUFX2 g_n677 (and_n291_n676, n677);
	INVX1 g_not_n1534 (n1534, not_n1534);
	BUFX2 g_n329 (and_n301_not_n328, n329);
	AND2X1 g_and_n379_not_n1082 (not_n1082, n379, and_n379_not_n1082);
	INVX1 g_not_n1325_3 (n1325, not_n1325_3);
	BUFX2 g_n1452 (and_not_pi065_0_not_pi138_6, n1452);
	AND2X1 g_and_not_n1500_not_n1501 (not_n1500, not_n1501, and_not_n1500_not_n1501);
	BUFX2 g_n408 (and_not_pi043_0_n407, n408);
	BUFX2 g_n1105 (and_not_pi024_4_not_pi042_2, n1105);
	BUFX2 g_n1146 (and_not_pi096_3_n1145, n1146);
	BUFX2 g_po125 (po125_driver, po125);
	INVX1 g_not_pi129_168830552257994114252669163302859949191483641195385604940410056010 (pi129, not_pi129_168830552257994114252669163302859949191483641195385604940410056010);
	INVX1 g_not_n1516 (n1516, not_n1516);
	BUFX2 g_n1148 (and_not_n1144_not_n1147, n1148);
	AND2X1 g_and_n390_n706 (n706, n390, and_n390_n706);
	INVX1 g_not_n1518 (n1518, not_n1518);
	BUFX2 g_n1399 (and_pi091_not_n1386_2, n1399);
	INVX1 g_not_pi129_26517308458596534717790233816010 (pi129, not_pi129_26517308458596534717790233816010);
	INVX1 g_not_n783 (n783, not_n783);
	BUFX2 g_n358 (and_pi005_not_n332, n358);
	BUFX2 g_po134_driver (and_not_pi129_57908879424491981188665523012880962572678888930017262494560649211430_not_n724, po134_driver);
	INVX1 g_not_pi024_0 (pi024, not_pi024_0);
	INVX1 g_not_n1544 (n1544, not_n1544);
	BUFX2 g_n791 (and_not_pi027_4_n737, n791);
	BUFX2 g_n1428 (and_pi096_not_n1423_0, n1428);
	AND2X1 g_and_not_pi012_2_n461 (n461, not_pi012_2, and_not_pi012_2_n461);
	BUFX2 g_n1261 (and_not_pi139_n1249, n1261);
	AND2X1 g_and_n638_n642 (n638, n642, and_n638_n642);
	BUFX2 g_n744 (and_not_n742_n743, n744);
	INVX1 g_not_n816 (n816, not_n816);
	INVX1 g_not_pi129_1299348114471230201171721456984490 (pi129, not_pi129_1299348114471230201171721456984490);
	INVX1 g_not_n1451 (n1451, not_n1451);
	BUFX2 g_n785 (and_not_pi129_332329305696010_not_n784, n785);
	AND2X1 g_and_not_pi056_0_not_n301 (not_n301, not_pi056_0, and_not_pi056_0_not_n301);
	INVX1 g_not_n511 (n511, not_n511);
	BUFX2 g_n1429 (and_pi146_n1414, n1429);
	INVX1 g_not_n1339 (n1339, not_n1339);
	AND2X1 g_and_not_n805_not_n806 (not_n806, not_n805, and_not_n805_not_n806);
	INVX1 g_not_n414 (n414, not_n414);
	AND2X1 g_and_pi014_not_pi054_9 (not_pi054_9, pi014, and_pi014_not_pi054_9);
	INVX1 g_not_n1490 (n1490, not_n1490);
	INVX1 g_not_n1067 (n1067, not_n1067);
	INVX1 g_not_pi040 (pi040, not_pi040);
	BUFX2 g_n1140 (and_pi052_not_n940_0, n1140);
	AND2X1 g_and_not_n933_n937 (not_n933, n937, and_not_n933_n937);
	AND2X1 g_and_pi011_not_pi054_6 (pi011, not_pi054_6, and_pi011_not_pi054_6);
	INVX1 g_not_pi054_24010 (pi054, not_pi054_24010);
	AND2X1 g_and_not_n1053_n1062 (not_n1053, n1062, and_not_n1053_n1062);
	BUFX2 g_n1009 (and_not_n379_7_not_n1008, n1009);
	AND2X1 g_and_not_n1231_not_n1232 (not_n1231, not_n1232, and_not_n1231_not_n1232);
	INVX1 g_not_pi129_492217353521848729599618551903381776068465426225614008572624070 (pi129, not_pi129_492217353521848729599618551903381776068465426225614008572624070);
	BUFX2 g_n330 (and_n300_n329, n330);
	INVX1 g_not_pi026_1 (pi026, not_pi026_1);
	AND2X1 g_and_n503_n513 (n513, n503, and_n503_n513);
	INVX1 g_not_pi106_4 (pi106, not_pi106_4);
	INVX1 g_not_pi106_0 (pi106, not_pi106_0);
	INVX1 g_not_pi006 (pi006, not_pi006);
	AND2X1 g_and_n934_n935 (n935, n934, and_n934_n935);
	BUFX2 g_po057_driver (and_not_n989_n998, po057_driver);
	INVX1 g_not_n1524 (n1524, not_n1524);
	INVX1 g_not_pi116_5 (pi116, not_pi116_5);
	AND2X1 g_and_not_pi003_332329305696010_n1373 (n1373, not_pi003_332329305696010, and_not_pi003_332329305696010_n1373);
	AND2X1 g_and_n389_n1012 (n389, n1012, and_n389_n1012);
	INVX1 g_not_n1050 (n1050, not_n1050);
	AND2X1 g_and_not_pi096_3_n1145 (not_pi096_3, n1145, and_not_pi096_3_n1145);
	BUFX2 g_n1522 (and_pi100_pi138, n1522);
	AND2X1 g_and_n479_n678 (n678, n479, and_n479_n678);
	BUFX2 g_n523 (and_pi011_not_pi054_6, n523);
	BUFX2 g_n832 (and_pi029_not_pi097_0, n832);
	INVX1 g_not_n1301 (n1301, not_n1301);
	AND2X1 g_and_not_pi058_3_not_n835 (not_n835, not_pi058_3, and_not_pi058_3_not_n835);
	AND2X1 g_and_n347_n417 (n417, n347, and_n347_n417);
	INVX1 g_not_pi116_0 (pi116, not_pi116_0);
	BUFX2 g_n434 (and_n356_n433, n434);
	INVX1 g_not_pi129_43181145673964365640352930977077280875522488490 (pi129, not_pi129_43181145673964365640352930977077280875522488490);
	BUFX2 g_n608 (and_n605_n607, n608);
	INVX1 g_not_pi019 (pi019, not_pi019);
	AND2X1 g_and_pi092_pi138 (pi138, pi092, and_pi092_pi138);
	BUFX2 g_n1477 (and_not_pi137_5_not_n1476, n1477);
	INVX1 g_not_n720 (n720, not_n720);
	INVX1 g_not_n836 (n836, not_n836);
	OR2X1 g_or_n1457_n1464 (n1464, n1457, or_n1457_n1464);
	INVX1 g_not_n940 (n940, not_n940);
	AND2X1 g_and_not_pi013_5_n450 (n450, not_pi013_5, and_not_pi013_5_n450);
	AND2X1 g_and_not_pi025_0_pi029 (pi029, not_pi025_0, and_not_pi025_0_pi029);
	INVX1 g_not_pi044_3 (pi044, not_pi044_3);
	INVX1 g_not_n1502 (n1502, not_n1502);
	AND2X1 g_and_n446_n453 (n453, n446, and_n446_n453);
	BUFX2 g_n472 (and_pi007_not_pi054_2, n472);
	BUFX2 g_n1476 (and_not_n1474_not_n1475, n1476);
	AND2X1 g_and_not_n379_70_not_n1070 (not_n1070, not_n379_70, and_not_n379_70_not_n1070);
	BUFX2 g_n1159 (and_not_n379_168070_not_n1158, n1159);
	INVX1 g_not_n1166 (n1166, not_n1166);
	BUFX2 g_n644 (and_n642_n643, n644);
	INVX1 g_not_n1020 (n1020, not_n1020);
	INVX1 g_not_pi136_10 (pi136, not_pi136_10);
	BUFX2 g_n858 (and_not_n854_not_n857, n858);
	AND2X1 g_and_not_pi129_332329305696010_not_n784 (not_pi129_332329305696010, not_n784, and_not_pi129_332329305696010_not_n784);
	BUFX2 g_n955 (and_n638_n954, n955);
	BUFX2 g_n302 (and_not_pi009_not_pi011, n302);
	BUFX2 g_po032_driver (and_not_pi003_70_n618, po032_driver);
	INVX1 g_not_pi022_1 (pi022, not_pi022_1);
	BUFX2 g_n480 (and_not_pi005_4_n479, n480);
	INVX1 g_not_pi129_11044276742439206463052992010 (pi129, not_pi129_11044276742439206463052992010);
	AND2X1 g_and_not_n897_not_n898 (not_n897, not_n898, and_not_n897_not_n898);
	INVX1 g_not_n1433 (n1433, not_n1433);
	BUFX2 g_n1101 (and_n705_n1100, n1101);
	AND2X1 g_and_not_n1545_not_n1546 (not_n1546, not_n1545, and_not_n1545_not_n1546);
	BUFX2 g_n342 (and_n311_n341, n342);
	BUFX2 g_n558 (and_not_pi016_1_n354, n558);
	INVX1 g_not_n1276 (n1276, not_n1276);
	AND2X1 g_and_not_pi038_not_pi050 (not_pi050, not_pi038, and_not_pi038_not_pi050);
	INVX1 g_not_n797 (n797, not_n797);
	INVX1 g_not_n1423_2 (n1423, not_n1423_2);
	BUFX2 g_po097_driver (and_not_pi129_881247870897231951843937366879128181133112010_not_n1344, po097_driver);
	BUFX2 g_n1091 (and_not_n379_490_not_n1090, n1091);
	BUFX2 g_po088_driver (or_pi129_n1306, po088_driver);
	INVX1 g_not_pi129_0 (pi129, not_pi129_0);
	BUFX2 g_n548 (and_not_pi025_0_pi029, n548);
	INVX1 g_not_n578 (n578, not_n578);
	BUFX2 g_n1527 (and_pi137_not_n1526, n1527);
	INVX1 g_not_n865 (n865, not_n865);
	INVX1 g_not_n1168 (n1168, not_n1168);
	AND2X1 g_and_not_pi010_1_n449 (not_pi010_1, n449, and_not_pi010_1_n449);
	INVX1 g_not_pi138_10 (pi138, not_pi138_10);
	AND2X1 g_and_pi026_n855 (n855, pi026, and_pi026_n855);
	OR2X1 g_or_pi003_not_n339 (not_n339, pi003, or_pi003_not_n339);
	AND2X1 g_and_not_pi095_not_pi100 (not_pi100, not_pi095, and_not_pi095_not_pi100);
	INVX1 g_not_n965 (n965, not_n965);
	BUFX2 g_n1015 (and_not_n1010_n1014, n1015);
	AND2X1 g_and_not_n357_not_n358 (not_n358, not_n357, and_not_n357_not_n358);
	BUFX2 g_n423 (and_n418_n422, n423);
	AND2X1 g_and_n611_n614 (n614, n611, and_n611_n614);
	INVX1 g_not_n1563 (n1563, not_n1563);
	BUFX2 g_po048 (po048_driver, po048);
	INVX1 g_not_pi058_10 (pi058, not_pi058_10);
	INVX1 g_not_n658 (n658, not_n658);
	AND2X1 g_and_pi082_not_n1030 (not_n1030, pi082, and_pi082_not_n1030);
	INVX1 g_not_pi070 (pi070, not_pi070);
	INVX1 g_not_pi073 (pi073, not_pi073);
	INVX1 g_not_pi007_4 (pi007, not_pi007_4);
	AND2X1 g_and_n408_n1001 (n408, n1001, and_n408_n1001);
	INVX1 g_not_n1392 (n1392, not_n1392);
	BUFX2 g_po071 (po071_driver, po071);
	BUFX2 g_n875 (and_pi099_pi106, n875);
	BUFX2 g_n717 (and_pi100_not_n716, n717);
	INVX1 g_not_n1167 (n1167, not_n1167);
	BUFX2 g_n1583 (and_pi082_n1582, n1583);
	AND2X1 g_and_n487_n493 (n493, n487, and_n487_n493);
	AND2X1 g_and_pi054_n300 (n300, pi054, and_pi054_n300);
	AND2X1 g_and_not_n1420_not_n1422 (not_n1420, not_n1422, and_not_n1420_not_n1422);
	AND2X1 g_and_pi025_not_pi116 (not_pi116, pi025, and_pi025_not_pi116);
	BUFX2 g_n1426 (and_not_n1424_not_n1425, n1426);
	AND2X1 g_and_not_n947_not_n951 (not_n947, not_n951, and_not_n947_not_n951);
	AND2X1 g_and_n737_n1207 (n737, n1207, and_n737_n1207);
	INVX1 g_not_n1590 (n1590, not_n1590);
	INVX1 g_not_n520 (n520, not_n520);
	INVX1 g_not_n1347 (n1347, not_n1347);
	BUFX2 g_n1497 (and_not_pi112_n1324, n1497);
	BUFX2 g_po017 (po017_driver, po017);
	INVX1 g_not_n468 (n468, not_n468);
	INVX1 g_not_n365 (n365, not_n365);
	AND2X1 g_and_n774_n1374 (n774, n1374, and_n774_n1374);
	INVX1 g_not_n1335 (n1335, not_n1335);
	AND2X1 g_and_not_pi047_1_n568 (not_pi047_1, n568, and_not_pi047_1_n568);
	INVX1 g_not_pi137_70 (pi137, not_pi137_70);
	AND2X1 g_and_n579_n919 (n919, n579, and_n579_n919);
	BUFX2 g_n1280 (and_pi068_not_n1247_3, n1280);
	INVX1 g_not_n835 (n835, not_n835);
	AND2X1 g_and_not_n672_not_n681 (not_n672, not_n681, and_not_n672_not_n681);
	INVX1 g_not_pi003_9 (pi003, not_pi003_9);
	BUFX2 g_n581 (and_n407_n580, n581);
	BUFX2 g_po114 (po114_driver, po114);
	BUFX2 g_n708 (and_n649_n707, n708);
	BUFX2 g_po072_driver (and_not_pi003_968890104070_n1203, po072_driver);
	BUFX2 g_n1142 (and_not_n1140_n1141, n1142);
	BUFX2 g_n1225 (and_n1223_n1224, n1225);
	BUFX2 g_po085_driver (or_pi129_n1293, po085_driver);
	BUFX2 g_n647 (and_not_n379_1_not_n646, n647);
	INVX1 g_not_pi129_3445521474652941107197329863323672432479257983579298060008368490 (pi129, not_pi129_3445521474652941107197329863323672432479257983579298060008368490);
	INVX1 g_not_pi129_1742514982336908143055105517947102601079450420187483430 (pi129, not_pi129_1742514982336908143055105517947102601079450420187483430);
	BUFX2 g_n910 (and_pi093_pi106, n910);
	AND2X1 g_and_pi082_not_n390 (pi082, not_n390, and_pi082_not_n390);
	INVX1 g_not_n646 (n646, not_n646);
	INVX1 g_not_n1454 (n1454, not_n1454);
	AND2X1 g_and_not_pi003_8_n555 (not_pi003_8, n555, and_not_pi003_8_n555);
	BUFX2 g_n462 (and_not_pi012_2_n461, n462);
	AND2X1 g_and_not_pi106_not_n863 (not_pi106, not_n863, and_not_pi106_not_n863);
	INVX1 g_not_n779 (n779, not_n779);
	AND2X1 g_and_pi068_not_n1247_3 (not_n1247_3, pi068, and_pi068_not_n1247_3);
	INVX1 g_not_n1247_1 (n1247, not_n1247_1);
	INVX1 g_not_n1065 (n1065, not_n1065);
	BUFX2 g_n392 (and_not_pi002_n391, n392);
	INVX1 g_not_pi116_1 (pi116, not_pi116_1);
	AND2X1 g_and_n447_n466 (n466, n447, and_n447_n466);
	AND2X1 g_and_pi058_pi116 (pi116, pi058, and_pi058_pi116);
	AND2X1 g_and_not_pi003_968890104070_n1203 (not_pi003_968890104070, n1203, and_not_pi003_968890104070_n1203);
	INVX1 g_not_n1557 (n1557, not_n1557);
	AND2X1 g_and_pi137_not_n1549 (pi137, not_n1549, and_pi137_not_n1549);
	BUFX2 g_n965 (and_pi082_not_n573, n965);
	BUFX2 g_n1300 (and_pi072_not_n1271_1, n1300);
	AND2X1 g_and_pi091_not_n1386_2 (not_n1386_2, pi091, and_pi091_not_n1386_2);
	AND2X1 g_and_not_n379_10_not_n1056 (not_n1056, not_n379_10, and_not_n379_10_not_n1056);
	INVX1 g_not_n1584 (n1584, not_n1584);
	INVX1 g_not_n379_5 (n379, not_n379_5);
	INVX1 g_not_pi138_4 (pi138, not_pi138_4);
	BUFX2 g_n1479 (and_not_pi138_8_not_n1478, n1479);
	AND2X1 g_and_not_pi136_168070_not_n1547 (not_pi136_168070, not_n1547, and_not_pi136_168070_not_n1547);
	AND2X1 g_and_not_pi053_3_not_n816 (not_n816, not_pi053_3, and_not_pi053_3_not_n816);
	AND2X1 g_and_n379_not_n693 (n379, not_n693, and_n379_not_n693);
	BUFX2 g_n976 (and_n403_n405, n976);
	INVX1 g_not_pi129_1435036016098684342856030763566710717400773837392460666392490 (pi129, not_pi129_1435036016098684342856030763566710717400773837392460666392490);
	BUFX2 g_po022 (po022_driver, po022);
	BUFX2 g_po055_driver (and_not_n953_n963, po055_driver);
	BUFX2 g_po049_driver (and_not_pi129_273687473400809163430_not_n894, po049_driver);
	BUFX2 g_n1525 (and_pi035_n1360, n1525);
	BUFX2 g_n486 (and_pi008_not_pi054_3, n486);
	AND2X1 g_and_pi007_not_pi054_2 (pi007, not_pi054_2, and_pi007_not_pi054_2);
	AND2X1 g_and_pi088_pi106 (pi088, pi106, and_pi088_pi106);
	INVX1 g_not_n1362 (n1362, not_n1362);
	BUFX2 g_n1351 (and_not_pi072_not_pi138_2, n1351);
	BUFX2 g_n1316 (and_pi076_not_n1271_5, n1316);
	BUFX2 g_n1600 (and_not_pi136_2824752490_pi140, n1600);
	BUFX2 g_n1192 (and_not_pi085_10_n1187, n1192);
	INVX1 g_not_n1208 (n1208, not_n1208);
	BUFX2 g_po024 (po024_driver, po024);
	AND2X1 g_and_not_n544_not_n553 (not_n544, not_n553, and_not_n544_not_n553);
	AND2X1 g_and_pi097_n1149 (n1149, pi097, and_pi097_n1149);
	AND2X1 g_and_n726_n787 (n726, n787, and_n726_n787);
	INVX1 g_not_n1222 (n1222, not_n1222);
	AND2X1 g_and_not_pi002_n391 (n391, not_pi002, and_not_pi002_n391);
	INVX1 g_not_n1386_3 (n1386, not_n1386_3);
	BUFX2 g_n993 (and_pi082_not_n992, n993);
	BUFX2 g_n1509 (and_not_pi138_10_not_n1508, n1509);
	AND2X1 g_and_not_pi045_4_not_n1033 (not_pi045_4, not_n1033, and_not_pi045_4_not_n1033);
	AND2X1 g_and_not_n753_not_n757 (not_n753, not_n757, and_not_n753_not_n757);
	BUFX2 g_n977 (and_pi041_pi082, n977);
	AND2X1 g_and_n1251_n1270 (n1251, n1270, and_n1251_n1270);
	INVX1 g_not_pi129_185621159210175743024531636712070 (pi129, not_pi129_185621159210175743024531636712070);
	AND2X1 g_and_not_pi071_0_not_pi138_24010 (not_pi138_24010, not_pi071_0, and_not_pi071_0_not_pi138_24010);
	BUFX2 g_po047_driver (and_not_pi129_5585458640832840070_not_n880, po047_driver);
	INVX1 g_not_n1421 (n1421, not_n1421);
	AND2X1 g_and_not_n794_0_not_n1570 (not_n794_0, not_n1570, and_not_n794_0_not_n1570);
	BUFX2 g_n824 (and_n743_n755, n824);
	AND2X1 g_and_pi143_n1414 (pi143, n1414, and_pi143_n1414);
	INVX1 g_not_n1620 (n1620, not_n1620);
	BUFX2 g_n1313 (and_not_pi144_0_n1271, n1313);
	AND2X1 g_and_pi043_n641 (n641, pi043, and_pi043_n641);
	BUFX2 g_n1539 (and_pi023_pi138, n1539);
	INVX1 g_not_pi012_5 (pi012, not_pi012_5);
	BUFX2 g_n802 (and_n776_n801, n802);
	INVX1 g_not_pi137_1 (pi137, not_pi137_1);
	INVX1 g_not_n822 (n822, not_n822);
	AND2X1 g_and_n416_n527 (n416, n527, and_n416_n527);
	AND2X1 g_and_pi059_not_pi116_70 (not_pi116_70, pi059, and_pi059_not_pi116_70);
	BUFX2 g_n487 (and_n369_n417, n487);
	BUFX2 g_n1620 (and_not_pi003_273687473400809163430_n1619, n1620);
	BUFX2 g_n1256 (and_not_pi142_n1249, n1256);
	AND2X1 g_and_pi090_not_n1386_1 (pi090, not_n1386_1, and_pi090_not_n1386_1);
	AND2X1 g_and_not_pi005_not_pi022 (not_pi005, not_pi022, and_not_pi005_not_pi022);
	BUFX2 g_n933 (and_pi074_n932, n933);
	INVX1 g_not_pi106 (pi106, not_pi106);
	BUFX2 g_n1629 (and_not_pi003_1915812313805664144010_not_n1628, n1629);
	AND2X1 g_and_not_n498_not_n507 (not_n507, not_n498, and_not_n498_not_n507);
	AND2X1 g_and_n398_n401 (n398, n401, and_n398_n401);
	AND2X1 g_and_not_pi129_4_not_n455 (not_n455, not_pi129_4, and_not_pi129_4_not_n455);
	AND2X1 g_and_not_pi003_2_n484 (not_pi003_2, n484, and_not_pi003_2_n484);
	INVX1 g_not_pi058_1 (pi058, not_pi058_1);
	BUFX2 g_n631 (and_not_pi019_1_n630, n631);
	AND2X1 g_and_pi082_not_pi137_3 (pi082, not_pi137_3, and_pi082_not_pi137_3);
	BUFX2 g_n882 (and_pi090_pi106, n882);
	BUFX2 g_n313 (and_n311_n312, n313);
	AND2X1 g_and_not_pi012_5_n606 (not_pi012_5, n606, and_not_pi012_5_n606);
	BUFX2 g_po066_driver (and_not_pi129_63668057609090279857414351392240010_not_n1138, po066_driver);
	INVX1 g_not_n1331 (n1331, not_n1331);
	AND2X1 g_and_n344_n561 (n344, n561, and_n344_n561);
	AND2X1 g_and_not_pi017_not_pi021 (not_pi021, not_pi017, and_not_pi017_not_pi021);
	BUFX2 g_n1233 (and_not_n1231_not_n1232, n1233);
	INVX1 g_not_n1343 (n1343, not_n1343);
	AND2X1 g_and_not_n1040_n1045 (n1045, not_n1040, and_not_n1040_n1045);
	AND2X1 g_and_pi122_pi127 (pi122, pi127, and_pi122_pi127);
	AND2X1 g_and_n526_n529 (n529, n526, and_n526_n529);
	AND2X1 g_and_pi028_not_pi116_3 (not_pi116_3, pi028, and_pi028_not_pi116_3);
	INVX1 g_not_n1152 (n1152, not_n1152);
	BUFX2 g_n725 (and_not_pi097_n724, n725);
	INVX1 g_not_n1125 (n1125, not_n1125);
	INVX1 g_not_pi140_0 (pi140, not_pi140_0);
	INVX1 g_not_n1442 (n1442, not_n1442);
	AND2X1 g_and_pi094_not_n1167 (pi094, not_n1167, and_pi094_not_n1167);
	BUFX2 g_n1490 (and_not_pi074_not_pi136_9, n1490);
	BUFX2 g_n431 (and_n416_n430, n431);
	INVX1 g_not_n1068 (n1068, not_n1068);
	BUFX2 g_po015_driver (or_pi003_not_n339, po015_driver);
	INVX1 g_not_pi011_4 (pi011, not_pi011_4);
	AND2X1 g_and_not_pi024_1_n380 (not_pi024_1, n380, and_not_pi024_1_n380);
	INVX1 g_not_n725 (n725, not_n725);
	BUFX2 g_n1210 (and_not_pi129_1070069044235980333563563003849377848070_not_n1209, n1210);
	BUFX2 g_po060_driver (and_not_n1034_n1046, po060_driver);
	AND2X1 g_and_not_pi003_47475615099430_n1234 (not_pi003_47475615099430, n1234, and_not_pi003_47475615099430_n1234);
	AND2X1 g_and_pi006_not_pi054_1 (pi006, not_pi054_1, and_pi006_not_pi054_1);
	INVX1 g_not_n1198 (n1198, not_n1198);
	BUFX2 g_n1170 (and_pi037_not_pi116_8, n1170);
	BUFX2 g_n296 (and_not_pi012_n295, n296);
	INVX1 g_not_pi085_7 (pi085, not_pi085_7);
	AND2X1 g_and_not_n657_not_n658 (not_n657, not_n658, and_not_n657_not_n658);
	BUFX2 g_n804 (and_not_n802_not_n803, n804);
	BUFX2 g_n978 (and_n390_n977, n978);
	INVX1 g_not_pi006_0 (pi006, not_pi006_0);
	BUFX2 g_po079 (po079_driver, po079);
	INVX1 g_not_n1271_1 (n1271, not_n1271_1);
	BUFX2 g_n306 (and_pi054_not_n305, n306);
	BUFX2 g_po050_driver (and_not_pi129_1915812313805664144010_not_n901, po050_driver);
	INVX1 g_not_n553 (n553, not_n553);
	INVX1 g_not_pi053_3 (pi053, not_pi053_3);
	INVX1 g_not_pi053_7 (pi053, not_pi053_7);
	BUFX2 g_n843 (and_pi053_not_pi058_4, n843);
	INVX1 g_not_pi068 (pi068, not_pi068);
	AND2X1 g_and_not_pi129_3119734822845423713013303218219760490_not_n1152 (not_n1152, not_pi129_3119734822845423713013303218219760490, and_not_pi129_3119734822845423713013303218219760490_not_n1152);
	AND2X1 g_and_pi100_pi138 (pi138, pi100, and_pi100_pi138);
	INVX1 g_not_n1386_0 (n1386, not_n1386_0);
	BUFX2 g_po065_driver (and_not_n1125_n1134, po065_driver);
	AND2X1 g_and_pi089_not_n1386_0 (not_n1386_0, pi089, and_pi089_not_n1386_0);
	BUFX2 g_po085 (po085_driver, po085);
	AND2X1 g_and_not_n1473_not_n1477 (not_n1477, not_n1473, and_not_n1473_not_n1477);
	AND2X1 g_and_pi063_n702 (pi063, n702, and_pi063_n702);
	INVX1 g_not_n896 (n896, not_n896);
	INVX1 g_not_n961 (n961, not_n961);
	AND2X1 g_and_not_pi136_57648010_pi139 (not_pi136_57648010, pi139, and_not_pi136_57648010_pi139);
	INVX1 g_not_n952 (n952, not_n952);
	AND2X1 g_and_pi111_not_n1421_0 (pi111, not_n1421_0, and_pi111_not_n1421_0);
	BUFX2 g_po048_driver (and_not_pi129_39098210485829880490_not_n887, po048_driver);
	INVX1 g_not_pi038_0 (pi038, not_pi038_0);
	BUFX2 g_po113 (po113_driver, po113);
	BUFX2 g_po071_driver (and_not_pi003_138412872010_n1185, po071_driver);
	INVX1 g_not_n846 (n846, not_n846);
	AND2X1 g_and_pi033_not_pi109_2 (pi033, not_pi109_2, and_pi033_not_pi109_2);
	AND2X1 g_and_n609_n615 (n615, n609, and_n609_n615);
	BUFX2 g_n433 (and_pi054_n300, n433);
	BUFX2 g_n1305 (and_not_pi141_0_n1271, n1305);
	AND2X1 g_and_not_n726_0_not_n792 (not_n726_0, not_n792, and_not_n726_0_not_n792);
	AND2X1 g_and_pi041_pi082 (pi041, pi082, and_pi041_pi082);
	AND2X1 g_and_n838_n843 (n838, n843, and_n838_n843);
	INVX1 g_not_n1010 (n1010, not_n1010);
	INVX1 g_not_n1022 (n1022, not_n1022);
	AND2X1 g_and_n390_n960 (n960, n390, and_n390_n960);
	INVX1 g_not_n334 (n334, not_n334);
	AND2X1 g_and_not_pi038_2_n641 (n641, not_pi038_2, and_not_pi038_2_n641);
	INVX1 g_not_pi129_21838143759917965991093122527538323430 (pi129, not_pi129_21838143759917965991093122527538323430);
	OR2X1 g_or_n1237_n1238 (n1238, n1237, or_n1237_n1238);
	INVX1 g_not_pi129_490 (pi129, not_pi129_490);
	AND2X1 g_and_pi069_not_n1247_4 (pi069, not_n1247_4, and_pi069_not_n1247_4);
	AND2X1 g_and_pi077_not_n1271_6 (not_n1271_6, pi077, and_pi077_not_n1271_6);
	AND2X1 g_and_not_pi144_0_n1271 (n1271, not_pi144_0, and_not_pi144_0_n1271);
	INVX1 g_not_pi129_29286449308136415160327158440136953416342323212091034008010 (pi129, not_pi129_29286449308136415160327158440136953416342323212091034008010);
	BUFX2 g_n1531 (and_not_n713_0_not_n1530, n1531);
	INVX1 g_not_pi129_63668057609090279857414351392240010 (pi129, not_pi129_63668057609090279857414351392240010);
	AND2X1 g_and_not_n1272_not_n1273 (not_n1273, not_n1272, and_not_n1272_not_n1273);
	INVX1 g_not_n1170 (n1170, not_n1170);
	BUFX2 g_po118_driver (or_n1484_n1494, po118_driver);
	BUFX2 g_n1219 (and_n726_n787, n1219);
	BUFX2 g_po023_driver (and_not_pi003_3_n496, po023_driver);
	BUFX2 g_n1485 (and_pi078_not_pi136_8, n1485);
	INVX1 g_not_pi054_5 (pi054, not_pi054_5);
	BUFX2 g_n353 (and_not_pi001_not_n352, n353);
	INVX1 g_not_n1463 (n1463, not_n1463);
	BUFX2 g_n985 (and_n927_n984, n985);
	BUFX2 g_po118 (po118_driver, po118);
	INVX1 g_not_n945 (n945, not_n945);
	BUFX2 g_po075 (po075_driver, po075);
	INVX1 g_not_pi129_2115876138024253916377293617876786762900601936010 (pi129, not_pi129_2115876138024253916377293617876786762900601936010);
	INVX1 g_not_n849 (n849, not_n849);
	INVX1 g_not_pi129_17984650426474121466202803405696493492512490 (pi129, not_pi129_17984650426474121466202803405696493492512490);
	AND2X1 g_and_pi000_not_pi123 (not_pi123, pi000, and_pi000_not_pi123);
	BUFX2 g_n535 (and_not_pi012_3_n449, n535);
	BUFX2 g_n525 (and_n448_n524, n525);
	BUFX2 g_n1361 (and_pi031_n1360, n1361);
	INVX1 g_not_pi013_3 (pi013, not_pi013_3);
	INVX1 g_not_n1109 (n1109, not_n1109);
	INVX1 g_not_pi106_9 (pi106, not_pi106_9);
	INVX1 g_not_n1325_5 (n1325, not_n1325_5);
	AND2X1 g_and_n499_n501 (n499, n501, and_n499_n501);
	INVX1 g_not_n1553 (n1553, not_n1553);
	AND2X1 g_and_not_pi009_2_n449 (n449, not_pi009_2, and_not_pi009_2_n449);
	AND2X1 g_and_not_pi024_3_n692 (not_pi024_3, n692, and_not_pi024_3_n692);
	BUFX2 g_n864 (and_not_pi106_not_n863, n864);
	BUFX2 g_n1512 (and_not_pi070_0_not_pi138_70, n1512);
	INVX1 g_not_pi054_490 (pi054, not_pi054_490);
	BUFX2 g_po031 (po031_driver, po031);
	INVX1 g_not_n695 (n695, not_n695);
	AND2X1 g_and_not_n595_not_n600 (not_n600, not_n595, and_not_n595_not_n600);
	AND2X1 g_and_pi119_pi138 (pi138, pi119, and_pi119_pi138);
	BUFX2 g_n1049 (and_n688_n927, n1049);
	BUFX2 g_n1628 (and_not_pi096_4_pi125, n1628);
	AND2X1 g_and_not_pi011_4_n418 (n418, not_pi011_4, and_not_pi011_4_n418);
	BUFX2 g_n816 (and_not_n809_not_n815, n816);
	AND2X1 g_and_not_pi129_1299348114471230201171721456984490_not_n1117 (not_pi129_1299348114471230201171721456984490, not_n1117, and_not_pi129_1299348114471230201171721456984490_not_n1117);
	INVX1 g_not_n913 (n913, not_n913);
	BUFX2 g_n1129 (and_not_n379_24010_not_n1128, n1129);
	BUFX2 g_n1516 (and_not_pi075_not_pi138_490, n1516);
	INVX1 g_not_n1613 (n1613, not_n1613);
	BUFX2 g_n335 (and_n302_not_n334, n335);
	BUFX2 g_po037 (po037_driver, po037);
	INVX1 g_not_n458 (n458, not_n458);
	INVX1 g_not_n1325 (n1325, not_n1325);
	AND2X1 g_and_pi076_not_n1271_5 (not_n1271_5, pi076, and_pi076_not_n1271_5);
	INVX1 g_not_pi022_3 (pi022, not_pi022_3);
	AND2X1 g_and_pi057_not_pi058_9 (pi057, not_pi058_9, and_pi057_not_pi058_9);
	AND2X1 g_and_pi027_pi116 (pi116, pi027, and_pi027_pi116);
	AND2X1 g_and_not_pi027_8_pi028 (not_pi027_8, pi028, and_not_pi027_8_pi028);
	BUFX2 g_n731 (and_pi026_n718, n731);
	BUFX2 g_n416 (and_not_pi009_1_not_pi014_3, n416);
	BUFX2 g_n737 (and_not_pi051_0_n736, n737);
	BUFX2 g_n1255 (and_pi063_not_n1247_0, n1255);
	INVX1 g_not_pi129_5 (pi129, not_pi129_5);
	AND2X1 g_and_not_n379_490_not_n1090 (not_n1090, not_n379_490, and_not_n379_490_not_n1090);
	INVX1 g_not_pi129_5080218607396233653221881976522165017724345248360010 (pi129, not_pi129_5080218607396233653221881976522165017724345248360010);
	AND2X1 g_and_not_pi006_not_pi007 (not_pi007, not_pi006, and_not_pi006_not_pi007);
	AND2X1 g_and_not_pi009_4_pi013 (pi013, not_pi009_4, and_not_pi009_4_pi013);
	INVX1 g_not_n893 (n893, not_n893);
	BUFX2 g_n1352 (and_not_n1350_not_n1351, n1352);
	BUFX2 g_po027 (po027_driver, po027);
	AND2X1 g_and_not_n1114_not_n1115 (not_n1115, not_n1114, and_not_n1114_not_n1115);
	INVX1 g_not_pi029 (pi029, not_pi029);
	AND2X1 g_and_not_pi129_21838143759917965991093122527538323430_not_n1184 (not_n1184, not_pi129_21838143759917965991093122527538323430, and_not_pi129_21838143759917965991093122527538323430_not_n1184);
	BUFX2 g_n484 (and_not_pi129_6_not_n483, n484);
	INVX1 g_not_pi077 (pi077, not_pi077);
	BUFX2 g_n899 (and_not_n897_not_n898, n899);
	INVX1 g_not_pi138_1176490 (pi138, not_pi138_1176490);
	BUFX2 g_po068_driver (and_not_pi026_10_n1155, po068_driver);
	INVX1 g_not_pi023 (pi023, not_pi023);
	BUFX2 g_n970 (and_n381_n405, n970);
	INVX1 g_not_pi137_4 (pi137, not_pi137_4);
	BUFX2 g_n1535 (and_not_pi071_0_not_pi138_24010, n1535);
	BUFX2 g_n1187 (and_not_pi026_3430_not_pi053_7, n1187);
	INVX1 g_not_n307 (n307, not_n307);
	INVX1 g_not_n1597 (n1597, not_n1597);
	INVX1 g_not_pi085_3 (pi085, not_pi085_3);
	AND2X1 g_and_pi050_n1041 (pi050, n1041, and_pi050_n1041);
	BUFX2 g_n1321 (and_not_pi146_0_n1271, n1321);
	BUFX2 g_po106_driver (and_not_pi129_5080218607396233653221881976522165017724345248360010_not_n1401, po106_driver);
	INVX1 g_not_n483 (n483, not_n483);
	AND2X1 g_and_not_pi003_168070_n683 (not_pi003_168070, n683, and_not_pi003_168070_n683);
	INVX1 g_not_n825 (n825, not_n825);
	AND2X1 g_and_not_pi129_43181145673964365640352930977077280875522488490_not_n1372 (not_n1372, not_pi129_43181145673964365640352930977077280875522488490, and_not_pi129_43181145673964365640352930977077280875522488490_not_n1372);
	INVX1 g_not_n1247 (n1247, not_n1247);
	INVX1 g_not_n1434 (n1434, not_n1434);
	BUFX2 g_n706 (and_pi024_pi082, n706);
	BUFX2 g_po028_driver (and_not_pi003_8_n555, po028_driver);
	BUFX2 g_n1117 (and_not_n1104_n1116, n1117);
	BUFX2 g_n311 (and_not_pi008_0_not_pi021_0, n311);
	INVX1 g_not_pi008_0 (pi008, not_pi008_0);
	AND2X1 g_and_n379_not_n921 (not_n921, n379, and_n379_not_n921);
	INVX1 g_not_n1500 (n1500, not_n1500);
	AND2X1 g_and_not_pi003_2326305139872070_not_n1246 (not_n1246, not_pi003_2326305139872070, and_not_pi003_2326305139872070_not_n1246);
	AND2X1 g_and_not_pi026_4_not_n723_0 (not_n723_0, not_pi026_4, and_not_pi026_4_not_n723_0);
	INVX1 g_not_n951 (n951, not_n951);
	INVX1 g_not_n1066 (n1066, not_n1066);
	INVX1 g_not_n1382 (n1382, not_n1382);
	INVX1 g_not_pi145 (pi145, not_pi145);
	INVX1 g_not_n1112 (n1112, not_n1112);
	INVX1 g_not_n1409 (n1409, not_n1409);
	INVX1 g_not_pi076 (pi076, not_pi076);
	INVX1 g_not_pi136_3 (pi136, not_pi136_3);
	BUFX2 g_n917 (and_pi082_not_n391, n917);
	INVX1 g_not_pi129_14811132966169777414641055325137507340304213552070 (pi129, not_pi129_14811132966169777414641055325137507340304213552070);
	INVX1 g_not_pi024_4 (pi024, not_pi024_4);
	AND2X1 g_and_not_pi129_302268019717750559482470516839540966128657419430_not_n1379 (not_pi129_302268019717750559482470516839540966128657419430, not_n1379, and_not_pi129_302268019717750559482470516839540966128657419430_not_n1379);
	AND2X1 g_and_not_pi017_0_n330 (not_pi017_0, n330, and_not_pi017_0_n330);
	INVX1 g_not_pi129_7490483309651862334944941026945644936490 (pi129, not_pi129_7490483309651862334944941026945644936490);
	BUFX2 g_n400 (and_n398_n399, n400);
	AND2X1 g_and_not_pi026_8_n749 (n749, not_pi026_8, and_not_pi026_8_n749);
	AND2X1 g_and_n418_n422 (n418, n422, and_n418_n422);
	INVX1 g_not_n700 (n700, not_n700);
	BUFX2 g_n1122 (and_pi082_not_n1121, n1122);
	INVX1 g_not_n1189 (n1189, not_n1189);
	INVX1 g_not_n1101 (n1101, not_n1101);
	AND2X1 g_and_n772_n774 (n772, n774, and_n772_n774);
	AND2X1 g_and_pi049_not_n1107 (not_n1107, pi049, and_pi049_not_n1107);
	BUFX2 g_n355 (and_not_pi008_1_not_pi011_1, n355);
	INVX1 g_not_n360 (n360, not_n360);
	BUFX2 g_n399 (and_not_pi047_0_not_pi048_0, n399);
	BUFX2 g_n1087 (and_n398_n401, n1087);
	BUFX2 g_n1359 (and_not_pi136_2_not_n1358, n1359);
	BUFX2 g_n584 (and_not_pi002_0_not_pi020_0, n584);
	BUFX2 g_n808 (and_not_n799_n807, n808);
	INVX1 g_not_n1305 (n1305, not_n1305);
	INVX1 g_not_pi129_3788186922656647816827176259430 (pi129, not_pi129_3788186922656647816827176259430);
	AND2X1 g_and_not_pi027_9_not_n845 (not_pi027_9, not_n845, and_not_pi027_9_not_n845);
	INVX1 g_not_n1031 (n1031, not_n1031);
	AND2X1 g_and_n302_not_n334 (n302, not_n334, and_n302_not_n334);
	AND2X1 g_and_not_n903_not_n907 (not_n903, not_n907, and_not_n903_not_n907);
	INVX1 g_not_n1330 (n1330, not_n1330);
	AND2X1 g_and_pi018_n295 (pi018, n295, and_pi018_n295);
	INVX1 g_not_pi129_39098210485829880490 (pi129, not_pi129_39098210485829880490);
	BUFX2 g_n596 (and_pi006_not_pi012_4, n596);
	AND2X1 g_and_pi037_not_pi116_8 (pi037, not_pi116_8, and_pi037_not_pi116_8);
	BUFX2 g_n1529 (and_n788_n1370, n1529);
	BUFX2 g_n871 (and_not_n869_not_n870, n871);
	BUFX2 g_n534 (and_pi012_not_pi054_7, n534);
	BUFX2 g_n1578 (and_not_pi003_797922662976120010_n1577, n1578);
	BUFX2 g_n762 (and_not_pi110_1_not_n761, n762);
	INVX1 g_not_pi047_2 (pi047, not_pi047_2);
	INVX1 g_not_pi116_6 (pi116, not_pi116_6);
	BUFX2 g_n662 (and_pi021_not_pi054_24010, n662);
	INVX1 g_not_n904 (n904, not_n904);
	INVX1 g_not_n1387 (n1387, not_n1387);
	INVX1 g_not_n371 (n371, not_n371);
	BUFX2 g_po138 (po138_driver, po138);
	AND2X1 g_and_not_pi053_not_n745 (not_pi053, not_n745, and_not_pi053_not_n745);
	BUFX2 g_n750 (and_not_pi027_0_n749, n750);
	INVX1 g_not_pi003_490 (pi003, not_pi003_490);
	AND2X1 g_and_pi120_pi138 (pi120, pi138, and_pi120_pi138);
	AND2X1 g_and_not_pi003_273687473400809163430_n1619 (n1619, not_pi003_273687473400809163430, and_not_pi003_273687473400809163430_n1619);
	INVX1 g_not_n1445 (n1445, not_n1445);
	AND2X1 g_and_not_pi064_not_pi138_8235430 (not_pi064, not_pi138_8235430, and_not_pi064_not_pi138_8235430);
	INVX1 g_not_n1142 (n1142, not_n1142);
	AND2X1 g_and_pi139_n1386 (pi139, n1386, and_pi139_n1386);
	BUFX2 g_n1317 (and_not_pi145_0_n1271, n1317);
	INVX1 g_not_n817 (n817, not_n817);
	BUFX2 g_n913 (and_not_n911_not_n912, n913);
	AND2X1 g_and_pi082_not_n1028 (not_n1028, pi082, and_pi082_not_n1028);
	AND2X1 g_and_pi035_pi109 (pi035, pi109, and_pi035_pi109);
	AND2X1 g_and_not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070_n1623 (n1623, not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070, and_not_pi129_2837535091800107078244610627631167166061265557570845862233471811360070_n1623);
	INVX1 g_not_n1416 (n1416, not_n1416);
	BUFX2 g_po036_driver (and_not_pi003_24010_n670, po036_driver);
	AND2X1 g_and_pi058_not_n839 (not_n839, pi058, and_pi058_not_n839);
	BUFX2 g_n1113 (and_not_n1108_not_n1112, n1113);
	INVX1 g_not_pi006_3 (pi006, not_pi006_3);
	INVX1 g_not_n957 (n957, not_n957);
	INVX1 g_not_n966 (n966, not_n966);
	AND2X1 g_and_not_pi050_4_not_n1124 (not_pi050_4, not_n1124, and_not_pi050_4_not_n1124);
	BUFX2 g_n690 (and_n573_n689, n690);
	AND2X1 g_and_not_pi096_4_pi125 (pi125, not_pi096_4, and_not_pi096_4_pi125);
	AND2X1 g_and_pi016_pi054 (pi016, pi054, and_pi016_pi054);
	BUFX2 g_po124_driver (and_pi116_n1573, po124_driver);
	BUFX2 g_n1374 (and_not_pi003_332329305696010_n1373, n1374);
	INVX1 g_not_n1422 (n1422, not_n1422);
	BUFX2 g_n473 (and_not_pi018_1_not_pi021_2, n473);
	INVX1 g_not_n408 (n408, not_n408);
	INVX1 g_not_pi137_5 (pi137, not_pi137_5);
	BUFX2 g_n705 (and_n583_n704, n705);
	INVX1 g_not_n1277 (n1277, not_n1277);
	AND2X1 g_and_pi034_pi136 (pi034, pi136, and_pi034_pi136);
	AND2X1 g_and_not_pi138_9_not_n1493 (not_pi138_9, not_n1493, and_not_pi138_9_not_n1493);
	INVX1 g_not_n1576 (n1576, not_n1576);
	INVX1 g_not_pi129_19773267430 (pi129, not_pi129_19773267430);
	BUFX2 g_n1011 (and_pi043_n641, n1011);
	INVX1 g_not_n1236 (n1236, not_n1236);
	BUFX2 g_po031_driver (and_not_pi003_10_n602, po031_driver);
	AND2X1 g_and_pi018_not_pi054_490 (not_pi054_490, pi018, and_pi018_not_pi054_490);
	BUFX2 g_n1249 (and_pi136_not_pi137_0, n1249);
	AND2X1 g_and_not_n1552_not_n1553 (not_n1552, not_n1553, and_not_n1552_not_n1553);
	BUFX2 g_n715 (and_not_pi096_n714, n715);
	BUFX2 g_n563 (and_n515_n562, n563);
	BUFX2 g_n914 (and_not_pi106_6_not_n913, n914);
	AND2X1 g_and_n478_n481 (n481, n478, and_n478_n481);
	INVX1 g_not_n1033 (n1033, not_n1033);
	AND2X1 g_and_n1246_not_n1591 (n1246, not_n1591, and_n1246_not_n1591);
	AND2X1 g_and_not_pi129_57648010_not_n635 (not_n635, not_pi129_57648010, and_not_pi129_57648010_not_n635);
	INVX1 g_not_pi054_4 (pi054, not_pi054_4);
	BUFX2 g_n793 (and_not_n726_0_not_n792, n793);
	INVX1 g_not_n1428 (n1428, not_n1428);
	AND2X1 g_and_not_pi129_9095436801298611408202050198891430_not_n1132 (not_n1132, not_pi129_9095436801298611408202050198891430, and_not_pi129_9095436801298611408202050198891430_not_n1132);
	AND2X1 g_and_pi116_not_n796_0 (pi116, not_n796_0, and_pi116_not_n796_0);
	AND2X1 g_and_not_n1191_not_n1193 (not_n1193, not_n1191, and_not_n1191_not_n1193);
	INVX1 g_not_pi071_0 (pi071, not_pi071_0);
	AND2X1 g_and_pi062_not_n1247 (pi062, not_n1247, and_pi062_not_n1247);
	BUFX2 g_n1102 (and_pi082_not_n1101, n1102);
	BUFX2 g_po133 (po133_driver, po133);
	BUFX2 g_n385 (and_n383_n384, n385);
	AND2X1 g_and_not_n989_n998 (n998, not_n989, and_not_n989_n998);
	BUFX2 g_n1588 (and_not_pi136_403536070_pi141, n1588);
	AND2X1 g_and_pi096_not_n1423_0 (pi096, not_n1423_0, and_pi096_not_n1423_0);
	BUFX2 g_n511 (and_pi010_not_pi054_5, n511);
	BUFX2 g_n1196 (and_pi060_n1144, n1196);
	AND2X1 g_and_not_pi050_1_n403 (not_pi050_1, n403, and_not_pi050_1_n403);
	BUFX2 g_po140_driver (and_not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430_not_n1629, po140_driver);
	AND2X1 g_and_pi005_not_pi007_9 (not_pi007_9, pi005, and_pi005_not_pi007_9);
	INVX1 g_not_pi050_0 (pi050, not_pi050_0);
	BUFX2 g_n749 (and_pi053_not_pi085_2, n749);
	AND2X1 g_and_not_n1444_not_n1445 (not_n1444, not_n1445, and_not_n1444_not_n1445);
	BUFX2 g_n1054 (and_not_pi050_3_n404, n1054);
	BUFX2 g_n820 (and_not_pi026_8_n749, n820);
	BUFX2 g_n848 (and_n787_n847, n848);
	AND2X1 g_and_n386_n393 (n386, n393, and_n386_n393);
	AND2X1 g_and_pi082_not_n948 (not_n948, pi082, and_pi082_not_n948);
	INVX1 g_not_n1477 (n1477, not_n1477);
	AND2X1 g_and_pi138_not_n1468 (pi138, not_n1468, and_pi138_not_n1468);
	AND2X1 g_and_pi084_not_pi136_70 (pi084, not_pi136_70, and_pi084_not_pi136_70);
	AND2X1 g_and_n1100_not_n1109 (not_n1109, n1100, and_n1100_not_n1109);
	BUFX2 g_n921 (and_pi082_not_n920, n921);
	INVX1 g_not_n379_168070 (n379, not_n379_168070);
	BUFX2 g_n1287 (and_n1251_n1286, n1287);
	AND2X1 g_and_not_n1377_not_n1378 (not_n1377, not_n1378, and_not_n1377_not_n1378);
	INVX1 g_not_pi065 (pi065, not_pi065);
	AND2X1 g_and_not_n1125_n1134 (not_n1125, n1134, and_not_n1125_n1134);
	AND2X1 g_and_not_n379_1_not_n646 (not_n646, not_n379_1, and_not_n379_1_not_n646);
	AND2X1 g_and_not_n1562_not_n1563 (not_n1562, not_n1563, and_not_n1562_not_n1563);
	BUFX2 g_n1466 (and_pi091_n1249, n1466);
	BUFX2 g_n580 (and_n570_n579, n580);
	AND2X1 g_and_not_po129_n1162 (n1162, not_po129, and_not_po129_n1162);
	INVX1 g_not_n1218 (n1218, not_n1218);
	INVX1 g_not_n1571 (n1571, not_n1571);
	AND2X1 g_and_n345_n597 (n597, n345, and_n345_n597);
	INVX1 g_not_pi038_2 (pi038, not_pi038_2);
	BUFX2 g_po135_driver (and_not_pi111_n1621, po135_driver);
	INVX1 g_not_pi142 (pi142, not_pi142);
	INVX1 g_not_pi110_1 (pi110, not_pi110_1);
	BUFX2 g_n928 (and_not_pi050_2_n391, n928);
	INVX1 g_not_n1309 (n1309, not_n1309);
	INVX1 g_not_n1537 (n1537, not_n1537);
	AND2X1 g_and_pi141_n1386 (n1386, pi141, and_pi141_n1386);
	INVX1 g_not_n541 (n541, not_n541);
	AND2X1 g_and_n445_n608 (n608, n445, and_n445_n608);
	AND2X1 g_and_not_n904_not_n905 (not_n905, not_n904, and_not_n904_not_n905);
	BUFX2 g_n1108 (and_pi049_not_n1107, n1108);
	AND2X1 g_and_n942_not_n944 (n942, not_n944, and_n942_not_n944);
	AND2X1 g_and_n345_n357 (n345, n357, and_n345_n357);
	BUFX2 g_n898 (and_pi035_not_pi109_4, n898);
	AND2X1 g_and_not_pi026_3_n787 (not_pi026_3, n787, and_not_pi026_3_n787);
	AND2X1 g_and_not_n310_not_n333 (not_n333, not_n310, and_not_n310_not_n333);
	AND2X1 g_and_not_pi136_24010_not_n1540 (not_pi136_24010, not_n1540, and_not_pi136_24010_not_n1540);
	INVX1 g_not_pi026_3 (pi026, not_pi026_3);
	BUFX2 g_n900 (and_not_pi106_4_not_n899, n900);
	AND2X1 g_and_not_n314_not_n315 (not_n314, not_n315, and_not_n314_not_n315);
	AND2X1 g_and_pi020_n411 (pi020, n411, and_pi020_n411);
	INVX1 g_not_pi085_10 (pi085, not_pi085_10);
	AND2X1 g_and_not_pi049_0_n383 (n383, not_pi049_0, and_not_pi049_0_n383);
	BUFX2 g_n1240 (and_not_pi114_pi123, n1240);
	BUFX2 g_n1309 (and_not_pi142_0_n1271, n1309);
	INVX1 g_not_n1504 (n1504, not_n1504);
	INVX1 g_not_pi061 (pi061, not_pi061);
	AND2X1 g_and_pi082_not_n1049 (pi082, not_n1049, and_pi082_not_n1049);
	BUFX2 g_n924 (and_not_pi038_1_not_n923, n924);
	AND2X1 g_and_pi025_not_pi029_0 (pi025, not_pi029_0, and_pi025_not_pi029_0);
	AND2X1 g_and_n406_n579 (n406, n579, and_n406_n579);
	INVX1 g_not_n889 (n889, not_n889);
	INVX1 g_not_n554 (n554, not_n554);
	INVX1 g_not_n1119 (n1119, not_n1119);
	INVX1 g_not_n1069 (n1069, not_n1069);
	BUFX2 g_n1557 (and_not_pi067_not_pi138_57648010, n1557);
	INVX1 g_not_n1547 (n1547, not_n1547);
	BUFX2 g_n401 (and_not_pi049_0_n383, n401);
	AND2X1 g_and_n432_n434 (n432, n434, and_n432_n434);
	AND2X1 g_and_pi060_not_n1236 (pi060, not_n1236, and_pi060_not_n1236);
	AND2X1 g_and_pi054_not_n305 (not_n305, pi054, and_pi054_not_n305);
	AND2X1 g_and_n612_n613 (n613, n612, and_n612_n613);
	AND2X1 g_and_n450_n621 (n450, n621, and_n450_n621);
	AND2X1 g_and_not_n313_not_n319 (not_n319, not_n313, and_not_n313_not_n319);
	AND2X1 g_and_n299_n665 (n299, n665, and_n299_n665);
	BUFX2 g_n572 (and_not_pi046_1_n388, n572);
	AND2X1 g_and_not_pi009_not_pi011 (not_pi011, not_pi009, and_not_pi009_not_pi011);
	AND2X1 g_and_not_pi039_0_not_pi052_0 (not_pi052_0, not_pi039_0, and_not_pi039_0_not_pi052_0);
	AND2X1 g_and_not_pi058_0_n773 (n773, not_pi058_0, and_not_pi058_0_n773);
	INVX1 g_not_n831 (n831, not_n831);
	BUFX2 g_n1164 (and_not_pi026_70_pi058, n1164);
	INVX1 g_not_n682 (n682, not_n682);
	AND2X1 g_and_n300_not_n371 (not_n371, n300, and_n300_not_n371);
	BUFX2 g_n842 (and_not_pi053_4_not_n841, n842);
	BUFX2 g_po105 (po105_driver, po105);
	AND2X1 g_and_not_pi106_7_not_n941 (not_pi106_7, not_n941, and_not_pi106_7_not_n941);
	BUFX2 g_n496 (and_not_pi129_7_not_n495, n496);
	AND2X1 g_and_n399_n704 (n704, n399, and_n399_n704);
	BUFX2 g_n1216 (and_not_n726_1_n787, n1216);
	INVX1 g_not_pi012 (pi012, not_pi012);
	AND2X1 g_and_not_pi038_1_not_n923 (not_pi038_1, not_n923, and_not_pi038_1_not_n923);
	BUFX2 g_n1051 (and_n379_not_n1050, n1051);
	BUFX2 g_po101_driver (and_not_pi129_302268019717750559482470516839540966128657419430_not_n1379, po101_driver);
	BUFX2 g_po096_driver (and_not_pi129_125892552985318850263419623839875454447587430_not_n1340, po096_driver);
	INVX1 g_not_n1608 (n1608, not_n1608);
	INVX1 g_not_pi129_2326305139872070 (pi129, not_pi129_2326305139872070);
	BUFX2 g_n1006 (and_not_pi047_2_n407, n1006);
	INVX1 g_not_pi027_5 (pi027, not_pi027_5);
	BUFX2 g_n904 (and_pi035_pi109, n904);
	BUFX2 g_po089_driver (or_pi129_n1310, po089_driver);
	BUFX2 g_n634 (and_n487_n633, n634);
	AND2X1 g_and_n388_n391 (n388, n391, and_n388_n391);
	AND2X1 g_and_not_n1524_not_n1525 (not_n1524, not_n1525, and_not_n1524_not_n1525);
	BUFX2 g_n1157 (and_n408_n1001, n1157);
	INVX1 g_not_pi138_5 (pi138, not_pi138_5);
	AND2X1 g_and_not_n1130_n1133 (not_n1130, n1133, and_not_n1130_n1133);
	AND2X1 g_and_not_pi106_2_not_n885 (not_n885, not_pi106_2, and_not_pi106_2_not_n885);
	AND2X1 g_and_pi015_not_n581 (not_n581, pi015, and_pi015_not_n581);
	BUFX2 g_n1226 (and_not_n1222_not_n1225, n1226);
	AND2X1 g_and_not_pi146_n1249 (n1249, not_pi146, and_not_pi146_n1249);
	BUFX2 g_n1183 (and_n1175_n1182, n1183);
	INVX1 g_not_n1491 (n1491, not_n1491);
	BUFX2 g_n740 (and_pi027_not_n739, n740);
	AND2X1 g_and_not_pi113_n426 (not_pi113, n426, and_not_pi113_n426);
	INVX1 g_not_n1313 (n1313, not_n1313);
	AND2X1 g_and_not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430_not_n1629 (not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430, not_n1629, and_not_pi129_139039219498205246833985920753927191137002012320971447249440118756643430_not_n1629);
	INVX1 g_not_pi058_3 (pi058, not_pi058_3);
	AND2X1 g_and_n934_n1011 (n1011, n934, and_n934_n1011);
	BUFX2 g_n557 (and_pi014_not_pi054_9, n557);
	BUFX2 g_n826 (and_not_n823_not_n825, n826);
	INVX1 g_not_n1567 (n1567, not_n1567);
	AND2X1 g_and_not_pi142_0_n1271 (n1271, not_pi142_0, and_not_pi142_0_n1271);
	BUFX2 g_n611 (and_n450_n610, n611);
	BUFX2 g_n1012 (and_n934_n1011, n1012);
	AND2X1 g_and_not_n307_not_n337 (not_n337, not_n307, and_not_n307_not_n337);
	AND2X1 g_and_not_n1451_not_n1455 (not_n1455, not_n1451, and_not_n1451_not_n1455);
	AND2X1 g_and_not_pi069_0_pi136 (not_pi069_0, pi136, and_not_pi069_0_pi136);
	BUFX2 g_po025 (po025_driver, po025);
	INVX1 g_not_pi012_1 (pi012, not_pi012_1);
	AND2X1 g_and_not_pi003_403536070_n827 (n827, not_pi003_403536070, and_not_pi003_403536070_n827);
	BUFX2 g_n1014 (and_not_pi129_11044276742439206463052992010_not_n1013, n1014);
	AND2X1 g_and_not_n397_not_n413 (not_n397, not_n413, and_not_n397_not_n413);
	BUFX2 g_n599 (and_n417_n598, n599);
	INVX1 g_not_n324 (n324, not_n324);
	AND2X1 g_and_pi036_not_pi109_5 (pi036, not_pi109_5, and_pi036_not_pi109_5);
	AND2X1 g_and_n459_n462 (n459, n462, and_n459_n462);
	AND2X1 g_and_not_n1589_not_n1590 (not_n1589, not_n1590, and_not_n1589_not_n1590);
	AND2X1 g_and_pi133_n1631 (n1631, pi133, and_pi133_n1631);
	AND2X1 g_and_pi082_not_n972 (pi082, not_n972, and_pi082_not_n972);
	INVX1 g_not_pi137_7 (pi137, not_pi137_7);
	BUFX2 g_n1045 (and_not_pi129_541169560379521116689596608490_not_n1044, n1045);
	BUFX2 g_n673 (and_not_pi022_3_n449, n673);
	INVX1 g_not_n887 (n887, not_n887);
	INVX1 g_not_pi024 (pi024, not_pi024);
	AND2X1 g_and_not_n728_0_n762 (n762, not_n728_0, and_not_n728_0_n762);
	AND2X1 g_and_pi095_not_pi096_1 (not_pi096_1, pi095, and_pi095_not_pi096_1);
	AND2X1 g_and_pi081_not_n1325_2 (not_n1325_2, pi081, and_pi081_not_n1325_2);
	BUFX2 g_n1346 (and_pi089_pi138, n1346);
	INVX1 g_not_n1448 (n1448, not_n1448);
	AND2X1 g_and_pi005_not_pi054_0 (pi005, not_pi054_0, and_pi005_not_pi054_0);
	INVX1 g_not_n379_7 (n379, not_n379_7);
	AND2X1 g_and_pi068_n1039 (n1039, pi068, and_pi068_n1039);
	BUFX2 g_po022_driver (and_not_pi003_2_n484, po022_driver);
	BUFX2 g_n1154 (and_not_pi003_19773267430_n1153, n1154);
	AND2X1 g_and_n416_n430 (n430, n416, and_n416_n430);
	BUFX2 g_n686 (and_not_pi129_138412872010_not_n685, n686);
	INVX1 g_not_n352 (n352, not_n352);
	AND2X1 g_and_not_n1521_not_n1522 (not_n1521, not_n1522, and_not_n1521_not_n1522);
	AND2X1 g_and_pi015_n411 (pi015, n411, and_pi015_n411);
	AND2X1 g_and_not_n1440_not_n1441 (not_n1440, not_n1441, and_not_n1440_not_n1441);
	BUFX2 g_n931 (and_pi082_not_n930, n931);
	AND2X1 g_and_not_n761_0_not_n1371 (not_n761_0, not_n1371, and_not_n761_0_not_n1371);
	AND2X1 g_and_not_pi136_2_not_n1358 (not_n1358, not_pi136_2, and_not_pi136_2_not_n1358);
	INVX1 g_not_n1440 (n1440, not_n1440);
	BUFX2 g_po141 (po141_driver, po141);
	INVX1 g_not_pi046 (pi046, not_pi046);
	BUFX2 g_n1291 (and_not_pi144_n1249, n1291);
	BUFX2 g_n1391 (and_pi089_not_n1386_0, n1391);
	AND2X1 g_and_pi139_n1325 (n1325, pi139, and_pi139_n1325);
	AND2X1 g_and_pi082_not_n1157 (pi082, not_n1157, and_pi082_not_n1157);
	AND2X1 g_and_not_pi046_2_not_n1052 (not_n1052, not_pi046_2, and_not_pi046_2_not_n1052);
	BUFX2 g_n589 (and_not_n582_not_n588, n589);
	AND2X1 g_and_not_pi019_1_n630 (n630, not_pi019_1, and_not_pi019_1_n630);
	INVX1 g_not_n1458 (n1458, not_n1458);
	AND2X1 g_and_not_pi129_1181813865805958799768684143120019644340385488367699234582870392070_not_n1608 (not_n1608, not_pi129_1181813865805958799768684143120019644340385488367699234582870392070, and_not_pi129_1181813865805958799768684143120019644340385488367699234582870392070_not_n1608);
	INVX1 g_not_pi046_0 (pi046, not_pi046_0);
	BUFX2 g_n398 (and_not_pi024_0_not_pi045_0, n398);
	AND2X1 g_and_n301_not_n302 (not_n302, n301, and_n301_not_n302);
	BUFX2 g_n716 (and_not_n713_not_n715, n716);
	AND2X1 g_and_pi085_not_n812 (pi085, not_n812, and_pi085_not_n812);
	INVX1 g_not_n620 (n620, not_n620);
	AND2X1 g_and_not_pi129_657123623635342801395430_not_n936 (not_pi129_657123623635342801395430, not_n936, and_not_pi129_657123623635342801395430_not_n936);
	BUFX2 g_n1404 (and_pi144_n1386, n1404);
	AND2X1 g_and_not_n410_not_n411 (not_n411, not_n410, and_not_n410_not_n411);
	INVX1 g_not_n839 (n839, not_n839);
	INVX1 g_not_pi129_597682638941559493067901192655856192170251494124306816490 (pi129, not_pi129_597682638941559493067901192655856192170251494124306816490);
	BUFX2 g_n412 (and_not_n410_not_n411, n412);
	INVX1 g_not_pi139_0 (pi139, not_pi139_0);
	BUFX2 g_n1519 (and_not_n1514_not_n1518, n1519);
	INVX1 g_not_n519 (n519, not_n519);
	INVX1 g_not_n1255 (n1255, not_n1255);
	INVX1 g_not_n1526 (n1526, not_n1526);
	AND2X1 g_and_not_n590_not_n591 (not_n591, not_n590, and_not_n590_not_n591);
	INVX1 g_not_n323 (n323, not_n323);
	AND2X1 g_and_not_pi013_0_not_n317 (not_pi013_0, not_n317, and_not_pi013_0_not_n317);
	INVX1 g_not_n654 (n654, not_n654);
	AND2X1 g_and_n1223_n1228 (n1223, n1228, and_n1223_n1228);
	INVX1 g_not_pi129_4183778472590916451475308348590993345191760458870147715430 (pi129, not_pi129_4183778472590916451475308348590993345191760458870147715430);
	AND2X1 g_and_pi025_not_pi026_1 (not_pi026_1, pi025, and_pi025_not_pi026_1);
	INVX1 g_not_n375 (n375, not_n375);
	AND2X1 g_and_not_n1092_n1097 (n1097, not_n1092, and_not_n1092_n1097);
	BUFX2 g_n1623 (and_pi081_pi120, n1623);
	BUFX2 g_n561 (and_not_pi009_4_pi013, n561);
	AND2X1 g_and_pi091_pi106 (pi106, pi091, and_pi091_pi106);
	INVX1 g_not_n1585 (n1585, not_n1585);
	INVX1 g_not_n864 (n864, not_n864);
	BUFX2 g_n1040 (and_pi068_n1039, n1040);
	INVX1 g_not_pi003_70 (pi003, not_pi003_70);
	INVX1 g_not_pi129_16284135979104490 (pi129, not_pi129_16284135979104490);
	BUFX2 g_n1366 (and_pi141_n1325, n1366);
	INVX1 g_not_n868 (n868, not_n868);
	AND2X1 g_and_n475_n477 (n477, n475, and_n475_n477);
	INVX1 g_not_pi129_9095436801298611408202050198891430 (pi129, not_pi129_9095436801298611408202050198891430);
	OR2X1 g_or_pi129_n1293 (pi129, n1293, or_pi129_n1293);
	BUFX2 g_n730 (and_not_n723_not_n729, n730);
	BUFX2 g_n478 (and_n475_n477, n478);
	INVX1 g_not_n995 (n995, not_n995);
	INVX1 g_not_pi042 (pi042, not_pi042);
	INVX1 g_not_n1386_2 (n1386, not_n1386_2);
	AND2X1 g_and_not_pi002_5_n383 (n383, not_pi002_5, and_not_pi002_5_n383);
	AND2X1 g_and_not_pi114_pi123 (pi123, not_pi114, and_not_pi114_pi123);
	BUFX2 g_n792 (and_not_n790_not_n791, n792);
	BUFX2 g_n906 (and_not_n904_not_n905, n906);
	INVX1 g_not_n1468 (n1468, not_n1468);
	AND2X1 g_and_not_pi138_10_not_n1508 (not_pi138_10, not_n1508, and_not_pi138_10_not_n1508);
	INVX1 g_not_n838 (n838, not_n838);
	BUFX2 g_n595 (and_pi016_not_pi054_10, n595);
	AND2X1 g_and_not_n1537_not_n1541 (not_n1537, not_n1541, and_not_n1537_not_n1541);
	BUFX2 g_n307 (and_not_pi000_not_n306, n307);
	INVX1 g_not_n1179 (n1179, not_n1179);
	INVX1 g_not_n1489 (n1489, not_n1489);
	INVX1 g_not_n379_2 (n379, not_n379_2);
	INVX1 g_not_pi129_403536070 (pi129, not_pi129_403536070);
	INVX1 g_not_pi001 (pi001, not_pi001);
	AND2X1 g_and_not_pi006_3_n341 (n341, not_pi006_3, and_not_pi006_3_n341);
	BUFX2 g_n1542 (and_not_n1537_not_n1541, n1542);
	INVX1 g_not_n1209 (n1209, not_n1209);
	BUFX2 g_po041 (po041_driver, po041);
	INVX1 g_not_n564 (n564, not_n564);
	BUFX2 g_n721 (and_not_pi026_not_n720, n721);
	BUFX2 g_n1288 (and_not_n1285_not_n1287, n1288);
	BUFX2 g_n1263 (and_not_n1260_not_n1262, n1263);
	AND2X1 g_and_pi085_not_pi116_1 (not_pi116_1, pi085, and_pi085_not_pi116_1);
	INVX1 g_not_n1601 (n1601, not_n1601);
	AND2X1 g_and_not_pi021_1_n300 (not_pi021_1, n300, and_not_pi021_1_n300);
	BUFX2 g_po123_driver (or_n1561_n1568, po123_driver);
	INVX1 g_not_pi141 (pi141, not_pi141);
	AND2X1 g_and_not_n1403_not_n1404 (not_n1404, not_n1403, and_not_n1403_not_n1404);
	INVX1 g_not_pi042_2 (pi042, not_pi042_2);
	AND2X1 g_and_pi017_n612 (pi017, n612, and_pi017_n612);
	AND2X1 g_and_not_pi069_n1103 (not_pi069, n1103, and_not_pi069_n1103);
	AND2X1 g_and_not_n379_24010_not_n1128 (not_n1128, not_n379_24010, and_not_n379_24010_not_n1128);
	INVX1 g_not_pi064 (pi064, not_pi064);
	INVX1 g_not_n616 (n616, not_n616);
	BUFX2 g_po064 (po064_driver, po064);
	AND2X1 g_and_not_pi026_10_n1155 (n1155, not_pi026_10, and_not_pi026_10_n1155);
	BUFX2 g_po009 (po009_driver, po009);
	AND2X1 g_and_n387_n388 (n388, n387, and_n387_n388);
	BUFX2 g_n795 (and_not_pi026_5_pi027, n795);
	AND2X1 g_and_not_pi116_4_n818 (n818, not_pi116_4, and_not_pi116_4_n818);
	AND2X1 g_and_pi019_n664 (n664, pi019, and_pi019_n664);
	BUFX2 g_po038_driver (and_pi061_n686, po038_driver);
	INVX1 g_not_pi010 (pi010, not_pi010);
	AND2X1 g_and_n298_n299 (n298, n299, and_n298_n299);
	AND2X1 g_and_not_n861_not_n862 (not_n862, not_n861, and_not_n861_not_n862);
	INVX1 g_not_pi044_1 (pi044, not_pi044_1);
	AND2X1 g_and_not_pi009_0_not_n367 (not_n367, not_pi009_0, and_not_pi009_0_not_n367);
	BUFX2 g_n1421 (and_pi138_n1412, n1421);
	AND2X1 g_and_pi030_n1360 (n1360, pi030, and_pi030_n1360);
	BUFX2 g_po013 (po013_driver, po013);
	BUFX2 g_po093 (po093_driver, po093);
	BUFX2 g_n1503 (and_not_pi137_7_not_n1502, n1503);
	BUFX2 g_po007 (po007_driver, po007);
	AND2X1 g_and_n448_n465 (n465, n448, and_n448_n465);
	AND2X1 g_and_not_pi129_492217353521848729599618551903381776068465426225614008572624070_n1586 (not_pi129_492217353521848729599618551903381776068465426225614008572624070, n1586, and_not_pi129_492217353521848729599618551903381776068465426225614008572624070_n1586);
	AND2X1 g_and_not_pi016_1_n354 (not_pi016_1, n354, and_not_pi016_1_n354);
	INVX1 g_not_pi046_2 (pi046, not_pi046_2);
	AND2X1 g_and_n503_n674 (n674, n503, and_n503_n674);
	AND2X1 g_and_n649_n707 (n707, n649, and_n649_n707);
	INVX1 g_not_n1381 (n1381, not_n1381);
	INVX1 g_not_n713_0 (n713, not_n713_0);
	BUFX2 g_n587 (and_n384_n586, n587);
	INVX1 g_not_n379_3 (n379, not_n379_3);
	AND2X1 g_and_pi052_not_n940_0 (not_n940_0, pi052, and_pi052_not_n940_0);
	AND2X1 g_and_pi132_pi133 (pi132, pi133, and_pi132_pi133);
	AND2X1 g_and_not_pi129_125892552985318850263419623839875454447587430_not_n1340 (not_n1340, not_pi129_125892552985318850263419623839875454447587430, and_not_pi129_125892552985318850263419623839875454447587430_not_n1340);
	AND2X1 g_and_pi090_n1249 (n1249, pi090, and_pi090_n1249);
	AND2X1 g_and_n447_n452 (n452, n447, and_n447_n452);
	AND2X1 g_and_n724_not_n833 (n724, not_n833, and_n724_not_n833);
	INVX1 g_not_pi136_6 (pi136, not_pi136_6);
	AND2X1 g_and_not_n1168_not_n1172 (not_n1168, not_n1172, and_not_n1168_not_n1172);
	BUFX2 g_n641 (and_not_pi040_1_not_pi042_0, n641);
	BUFX2 g_n1526 (and_not_n1524_not_n1525, n1526);
	AND2X1 g_and_not_pi029_1_pi059 (pi059, not_pi029_1, and_not_pi029_1_pi059);
	BUFX2 g_po088 (po088_driver, po088);
	INVX1 g_not_pi028_1 (pi028, not_pi028_1);
	INVX1 g_not_pi065_0 (pi065, not_pi065_0);
	INVX1 g_not_n1496 (n1496, not_n1496);
	INVX1 g_not_n435 (n435, not_n435);
	BUFX2 g_n1195 (and_pi057_not_n1194, n1195);
	INVX1 g_not_pi048 (pi048, not_pi048);
	BUFX2 g_n1363 (and_pi137_not_n1362, n1363);
	BUFX2 g_n813 (and_pi085_not_n812, n813);
	AND2X1 g_and_not_n1387_not_n1388 (not_n1387, not_n1388, and_not_n1387_not_n1388);
	AND2X1 g_and_not_n379_7_not_n1008 (not_n1008, not_n379_7, and_not_n379_7_not_n1008);
	AND2X1 g_and_not_pi137_4_not_n1456 (not_n1456, not_pi137_4, and_not_pi137_4_not_n1456);
	AND2X1 g_and_n514_n518 (n514, n518, and_n514_n518);
	AND2X1 g_and_not_n1304_not_n1305 (not_n1304, not_n1305, and_not_n1304_not_n1305);
	AND2X1 g_and_n459_n479 (n459, n479, and_n459_n479);
	INVX1 g_not_n1151 (n1151, not_n1151);
	AND2X1 g_and_pi073_not_n1271_2 (not_n1271_2, pi073, and_pi073_not_n1271_2);
	INVX1 g_not_n350 (n350, not_n350);
	AND2X1 g_and_not_n1365_not_n1366 (not_n1366, not_n1365, and_not_n1365_not_n1366);
	INVX1 g_not_n956 (n956, not_n956);
	INVX1 g_not_n1193 (n1193, not_n1193);
	AND2X1 g_and_n638_n1027 (n638, n1027, and_n638_n1027);
	AND2X1 g_and_not_n1346_not_n1347 (not_n1346, not_n1347, and_not_n1346_not_n1347);
	INVX1 g_not_pi053_8 (pi053, not_pi053_8);
	BUFX2 g_n1548 (and_not_pi136_168070_not_n1547, n1548);
	AND2X1 g_and_pi082_not_n700 (not_n700, pi082, and_pi082_not_n700);
	AND2X1 g_and_pi136_not_n1554 (pi136, not_n1554, and_pi136_not_n1554);
	BUFX2 g_n1448 (and_pi124_pi138, n1448);
	INVX1 g_not_pi129_332329305696010 (pi129, not_pi129_332329305696010);
	BUFX2 g_n1532 (and_not_pi129_1435036016098684342856030763566710717400773837392460666392490_not_n1531, n1532);
	BUFX2 g_n1621 (and_not_pi129_405362155971443868320658661090166738008752222510120837461924544480010_not_n1620, n1621);
	INVX1 g_not_n1205 (n1205, not_n1205);
	INVX1 g_not_pi009_3 (pi009, not_pi009_3);
	INVX1 g_not_pi106_7 (pi106, not_pi106_7);
	AND2X1 g_and_n389_n392 (n389, n392, and_n389_n392);
	INVX1 g_not_n1028 (n1028, not_n1028);
	AND2X1 g_and_not_n842_not_n844 (not_n844, not_n842, and_not_n842_not_n844);
	BUFX2 g_n709 (and_n705_n708, n709);
	AND2X1 g_and_pi027_n838 (n838, pi027, and_pi027_n838);
	BUFX2 g_po131_driver (and_pi054_n1610, po131_driver);
	BUFX2 g_n886 (and_not_pi106_2_not_n885, n886);
	BUFX2 g_n1232 (and_n856_n1223, n1232);
	AND2X1 g_and_not_pi048_1_n381 (not_pi048_1, n381, and_not_pi048_1_n381);
	AND2X1 g_and_not_n379_3_not_n931 (not_n931, not_n379_3, and_not_n379_3_not_n931);
	INVX1 g_not_n767 (n767, not_n767);
	BUFX2 g_po132_driver (or_not_pi122_2_pi129, po132_driver);
	AND2X1 g_and_pi060_n1144 (n1144, pi060, and_pi060_n1144);
	AND2X1 g_and_not_pi026_7_not_pi027_7 (not_pi026_7, not_pi027_7, and_not_pi026_7_not_pi027_7);
	AND2X1 g_and_not_pi005_3_not_pi007_5 (not_pi007_5, not_pi005_3, and_not_pi005_3_not_pi007_5);
	INVX1 g_not_pi017_0 (pi017, not_pi017_0);
	INVX1 g_not_pi041_2 (pi041, not_pi041_2);
	AND2X1 g_and_pi082_not_n1037 (pi082, not_n1037, and_pi082_not_n1037);
	INVX1 g_not_n305 (n305, not_n305);
	BUFX2 g_n1077 (and_not_pi129_26517308458596534717790233816010_not_n1076, n1077);
	AND2X1 g_and_n356_n433 (n433, n356, and_n356_n433);
	INVX1 g_not_n325 (n325, not_n325);
	INVX1 g_not_n366 (n366, not_n366);
	AND2X1 g_and_n400_n401 (n400, n401, and_n400_n401);
	BUFX2 g_n437 (and_not_n435_not_n436, n437);
	BUFX2 g_n1130 (and_pi066_n1129, n1130);
	AND2X1 g_and_n1251_n1261 (n1251, n1261, and_n1251_n1261);
	BUFX2 g_n1534 (and_pi098_pi138, n1534);
	INVX1 g_not_n1628 (n1628, not_n1628);
	BUFX2 g_po000 (po000_driver, po000);
	BUFX2 g_po069_driver (or_pi129_n1159, po069_driver);
	BUFX2 g_n1013 (and_n389_n1012, n1013);
	BUFX2 g_po017_driver (and_not_pi129_1_not_n414, po017_driver);
	BUFX2 g_n1546 (and_pi097_pi138, n1546);
	INVX1 g_not_pi058_8 (pi058, not_pi058_8);
	BUFX2 g_n1308 (and_pi074_not_n1271_3, n1308);
	INVX1 g_not_pi022_0 (pi022, not_pi022_0);
	INVX1 g_not_n744 (n744, not_n744);
	AND2X1 g_and_pi100_not_n1423_2 (not_n1423_2, pi100, and_pi100_not_n1423_2);
	BUFX2 g_po130_driver (and_not_pi129_168830552257994114252669163302859949191483641195385604940410056010_n1604, po130_driver);
	AND2X1 g_and_not_pi014_0_not_n320 (not_pi014_0, not_n320, and_not_pi014_0_not_n320);
	INVX1 g_not_n1325_6 (n1325, not_n1325_6);
	BUFX2 g_n872 (and_not_pi106_0_not_n871, n872);
	INVX1 g_not_n784 (n784, not_n784);
	BUFX2 g_n600 (and_n434_n599, n600);
	AND2X1 g_and_not_pi129_93874803376477543056490_not_n915 (not_pi129_93874803376477543056490, not_n915, and_not_pi129_93874803376477543056490_not_n915);
	INVX1 g_not_pi027_6 (pi027, not_pi027_6);
	INVX1 g_not_pi003_113988951853731430 (pi003, not_pi003_113988951853731430);
	INVX1 g_not_n1575 (n1575, not_n1575);
	INVX1 g_not_n691 (n691, not_n691);
	INVX1 g_not_n936 (n936, not_n936);
	INVX1 g_not_pi002_5 (pi002, not_pi002_5);
	INVX1 g_not_n944 (n944, not_n944);
	INVX1 g_not_n1199 (n1199, not_n1199);
	BUFX2 g_n529 (and_n369_n528, n529);
	INVX1 g_not_pi054_1 (pi054, not_pi054_1);
	AND2X1 g_and_n487_n633 (n487, n633, and_n487_n633);
	BUFX2 g_n803 (and_n728_n737, n803);
	BUFX2 g_n524 (and_not_pi011_3_n449, n524);
	INVX1 g_not_n854 (n854, not_n854);
	INVX1 g_not_n672 (n672, not_n672);
	BUFX2 g_po116_driver (or_n1457_n1464, po116_driver);
	AND2X1 g_and_not_n917_not_n922 (not_n922, not_n917, and_not_n917_not_n922);
	INVX1 g_not_pi143 (pi143, not_pi143);
	INVX1 g_not_n877 (n877, not_n877);
	AND2X1 g_and_pi144_n1414 (n1414, pi144, and_pi144_n1414);
	INVX1 g_not_n1312 (n1312, not_n1312);
	INVX1 g_not_pi003_10 (pi003, not_pi003_10);
	INVX1 g_not_n790 (n790, not_n790);
	AND2X1 g_and_pi010_not_pi022_1 (pi010, not_pi022_1, and_pi010_not_pi022_1);
	BUFX2 g_n300 (and_n298_n299, n300);
	AND2X1 g_and_n449_n558 (n558, n449, and_n449_n558);
	AND2X1 g_and_n300_n329 (n329, n300, and_n300_n329);
	AND2X1 g_and_not_pi013_4_n417 (n417, not_pi013_4, and_not_pi013_4_n417);
	AND2X1 g_and_pi051_not_pi109_7 (pi051, not_pi109_7, and_pi051_not_pi109_7);
	BUFX2 g_n1055 (and_n1049_n1054, n1055);
	AND2X1 g_and_pi080_not_n1325_1 (pi080, not_n1325_1, and_pi080_not_n1325_1);
	AND2X1 g_and_not_pi058_not_n752 (not_n752, not_pi058, and_not_pi058_not_n752);
	AND2X1 g_and_not_pi015_2_not_pi049_1 (not_pi049_1, not_pi015_2, and_not_pi015_2_not_pi049_1);
	INVX1 g_not_n769 (n769, not_n769);
	BUFX2 g_po052 (po052_driver, po052);
	INVX1 g_not_n1201 (n1201, not_n1201);
	AND2X1 g_and_n434_n599 (n434, n599, and_n434_n599);
	INVX1 g_not_n692 (n692, not_n692);
	AND2X1 g_and_not_n458_not_n468 (not_n468, not_n458, and_not_n458_not_n468);
	BUFX2 g_po016_driver (or_pi003_not_n377, po016_driver);
	INVX1 g_not_n379_1 (n379, not_n379_1);
	BUFX2 g_n884 (and_pi033_not_pi109_2, n884);
	BUFX2 g_n554 (and_not_n544_not_n553, n554);
	AND2X1 g_and_pi039_not_n943 (not_n943, pi039, and_pi039_not_n943);
	BUFX2 g_po097 (po097_driver, po097);
	BUFX2 g_n547 (and_n447_n546, n547);
	BUFX2 g_n1038 (and_pi082_not_n1037, n1038);
	AND2X1 g_and_n398_n925 (n925, n398, and_n398_n925);
	INVX1 g_not_pi138_3 (pi138, not_pi138_3);
	INVX1 g_not_pi136_70 (pi136, not_pi136_70);
	BUFX2 g_n972 (and_n927_n971, n972);
	INVX1 g_not_n734 (n734, not_n734);
	BUFX2 g_n812 (and_not_n810_not_n811, n812);
	INVX1 g_not_n953 (n953, not_n953);
	BUFX2 g_n463 (and_n459_n462, n463);
	BUFX2 g_n1082 (and_pi082_not_n919, n1082);
	BUFX2 g_n629 (and_pi017_n612, n629);
	AND2X1 g_and_not_pi129_47475615099430_not_n770 (not_pi129_47475615099430, not_n770, and_not_pi129_47475615099430_not_n770);
	INVX1 g_not_pi016 (pi016, not_pi016);
	BUFX2 g_n1434 (and_not_n1432_not_n1433, n1434);
	BUFX2 g_n1162 (and_pi114_not_pi122, n1162);
	INVX1 g_not_n1429 (n1429, not_n1429);
	INVX1 g_not_pi116_9 (pi116, not_pi116_9);
	BUFX2 g_n1178 (and_not_pi085_7_not_n1177, n1178);
	INVX1 g_not_n1252 (n1252, not_n1252);
	AND2X1 g_and_not_pi007_1_n311 (n311, not_pi007_1, and_not_pi007_1_n311);
	BUFX2 g_n1499 (and_pi138_not_n1498, n1499);
	BUFX2 g_po067_driver (and_not_pi129_445676403263631959001900459745680070_not_n1142, po067_driver);
	AND2X1 g_and_pi082_not_n1018 (not_n1018, pi082, and_pi082_not_n1018);
	BUFX2 g_n1563 (and_pi111_pi138, n1563);
	INVX1 g_not_pi017_4 (pi017, not_pi017_4);
	INVX1 g_not_pi122_0 (pi122, not_pi122_0);
	AND2X1 g_and_not_n746_not_n751 (not_n751, not_n746, and_not_n746_not_n751);
	BUFX2 g_n1100 (and_n384_n1054, n1100);
	AND2X1 g_and_pi026_n768 (n768, pi026, and_pi026_n768);
	INVX1 g_not_pi129_3119734822845423713013303218219760490 (pi129, not_pi129_3119734822845423713013303218219760490);
	INVX1 g_not_pi138_403536070 (pi138, not_pi138_403536070);
	BUFX2 g_po014 (po014_driver, po014);
	AND2X1 g_and_n787_n1175 (n787, n1175, and_n787_n1175);
	AND2X1 g_and_pi099_n1249 (n1249, pi099, and_pi099_n1249);
	INVX1 g_not_pi058_2 (pi058, not_pi058_2);
	AND2X1 g_and_not_n817_not_n821 (not_n821, not_n817, and_not_n817_not_n821);
	INVX1 g_not_n412 (n412, not_n412);
	AND2X1 g_and_not_n802_not_n803 (not_n803, not_n802, and_not_n802_not_n803);
	BUFX2 g_po125_driver (and_pi116_n1578, po125_driver);
	INVX1 g_not_n1034 (n1034, not_n1034);
	BUFX2 g_n1405 (and_not_n1403_not_n1404, n1405);
	BUFX2 g_n1412 (and_not_pi136_3_n1411, n1412);
	AND2X1 g_and_not_pi056_n308 (n308, not_pi056, and_not_pi056_n308);
	INVX1 g_not_pi003_6 (pi003, not_pi003_6);
	INVX1 g_not_n1535 (n1535, not_n1535);
	BUFX2 g_n498 (and_pi009_not_pi054_4, n498);
	AND2X1 g_and_not_pi073_not_pi136_10 (not_pi136_10, not_pi073, and_not_pi073_not_pi136_10);
	BUFX2 g_po087 (po087_driver, po087);
	BUFX2 g_n438 (and_not_pi129_3_not_n437, n438);
	BUFX2 g_n897 (and_pi034_pi109, n897);
	INVX1 g_not_n1386_5 (n1386, not_n1386_5);
	AND2X1 g_and_not_pi143_n1271 (not_pi143, n1271, and_not_pi143_n1271);
	BUFX2 g_n468 (and_n464_n467, n468);
	INVX1 g_not_pi114 (pi114, not_pi114);
	BUFX2 g_po105_driver (and_not_pi129_725745515342319093317411710931737859674906464051430_not_n1397, po105_driver);
	INVX1 g_not_pi136_4 (pi136, not_pi136_4);
	BUFX2 g_n552 (and_n550_n551, n552);
	INVX1 g_not_n1247_5 (n1247, not_n1247_5);
	INVX1 g_not_pi011_1 (pi011, not_pi011_1);
	INVX1 g_not_n920 (n920, not_n920);
	BUFX2 g_n1007 (and_n927_n1006, n1007);
	BUFX2 g_n1270 (and_not_pi136_not_pi137_1, n1270);
	INVX1 g_not_pi137_2 (pi137, not_pi137_2);
	OR2X1 g_or_pi129_n1268 (pi129, n1268, or_pi129_n1268);
	INVX1 g_not_n1247_0 (n1247, not_n1247_0);
	BUFX2 g_po095 (po095_driver, po095);
	BUFX2 g_po121_driver (and_not_pi003_16284135979104490_n1532, po121_driver);
	INVX1 g_not_n1393 (n1393, not_n1393);
	INVX1 g_not_pi005_1 (pi005, not_pi005_1);
	BUFX2 g_po009_driver (pi121, po009_driver);
	INVX1 g_not_pi040_1 (pi040, not_pi040_1);
	BUFX2 g_n958 (and_not_n379_4_not_n957, n958);
	BUFX2 g_n1419 (and_not_pi003_2326305139872070_not_n1246, n1419);
	BUFX2 g_po109 (po109_driver, po109);
	AND2X1 g_and_not_pi129_205005145156954906122290109080958673914396262484637238056070_not_n1446 (not_n1446, not_pi129_205005145156954906122290109080958673914396262484637238056070, and_not_pi129_205005145156954906122290109080958673914396262484637238056070_not_n1446);
	AND2X1 g_and_not_pi054_8235430_pi118 (not_pi054_8235430, pi118, and_not_pi054_8235430_pi118);
	BUFX2 g_n515 (and_n459_n479, n515);
	INVX1 g_not_pi009_2 (pi009, not_pi009_2);
	BUFX2 g_n582 (and_pi015_not_n581, n582);
	INVX1 g_not_n1357 (n1357, not_n1357);
	AND2X1 g_and_not_n1466_not_n1467 (not_n1466, not_n1467, and_not_n1466_not_n1467);
	BUFX2 g_n1590 (and_not_pi112_0_not_n1421_1, n1590);
	INVX1 g_not_pi003_1915812313805664144010 (pi003, not_pi003_1915812313805664144010);
	BUFX2 g_n984 (and_n688_n976, n984);
	BUFX2 g_n700 (and_n408_n699, n700);
	AND2X1 g_and_not_pi129_1_not_n414 (not_pi129_1, not_n414, and_not_pi129_1_not_n414);
	AND2X1 g_and_not_pi129_881247870897231951843937366879128181133112010_not_n1344 (not_n1344, not_pi129_881247870897231951843937366879128181133112010, and_not_pi129_881247870897231951843937366879128181133112010_not_n1344);
	AND2X1 g_and_not_n723_not_n729 (not_n723, not_n729, and_not_n723_not_n729);
	INVX1 g_not_pi025_0 (pi025, not_pi025_0);
	BUFX2 g_po008_driver (pi126, po008_driver);
	AND2X1 g_and_not_pi007_8_n346 (n346, not_pi007_8, and_not_pi007_8_n346);
	INVX1 g_not_n1326 (n1326, not_n1326);
	AND2X1 g_and_n447_n546 (n546, n447, and_n447_n546);
	BUFX2 g_n428 (and_not_n425_not_n427, n428);
	BUFX2 g_n1295 (and_pi071_not_n1247_6, n1295);
	AND2X1 g_and_not_pi137_5_not_n1476 (not_n1476, not_pi137_5, and_not_pi137_5_not_n1476);
	AND2X1 g_and_not_pi129_63668057609090279857414351392240010_not_n1138 (not_n1138, not_pi129_63668057609090279857414351392240010, and_not_pi129_63668057609090279857414351392240010_not_n1138);
	INVX1 g_not_n872 (n872, not_n872);
	AND2X1 g_and_not_pi129_17984650426474121466202803405696493492512490_not_n1336 (not_n1336, not_pi129_17984650426474121466202803405696493492512490, and_not_pi129_17984650426474121466202803405696493492512490_not_n1336);
	BUFX2 g_po121 (po121_driver, po121);
	AND2X1 g_and_pi082_not_n1007 (pi082, not_n1007, and_pi082_not_n1007);
	INVX1 g_not_n1399 (n1399, not_n1399);
	INVX1 g_not_n1415 (n1415, not_n1415);
	AND2X1 g_and_not_pi129_5080218607396233653221881976522165017724345248360010_not_n1401 (not_n1401, not_pi129_5080218607396233653221881976522165017724345248360010, and_not_pi129_5080218607396233653221881976522165017724345248360010_not_n1401);
	INVX1 g_not_n931 (n931, not_n931);
	BUFX2 g_po046 (po046_driver, po046);
	AND2X1 g_and_not_n1407_not_n1408 (not_n1408, not_n1407, and_not_n1407_not_n1408);
	INVX1 g_not_pi015_0 (pi015, not_pi015_0);
	AND2X1 g_and_not_pi129_24010_not_n593 (not_pi129_24010, not_n593, and_not_pi129_24010_not_n593);
	INVX1 g_not_pi129_12197604876358357001385738625629718207556152941312384010 (pi129, not_pi129_12197604876358357001385738625629718207556152941312384010);
	BUFX2 g_po051 (po051_driver, po051);
	BUFX2 g_po136 (po136_driver, po136);
	AND2X1 g_and_not_pi100_0_not_n781 (not_n781, not_pi100_0, and_not_pi100_0_not_n781);
	AND2X1 g_and_n408_n1036 (n1036, n408, and_n408_n1036);
	BUFX2 g_po025_driver (and_not_pi003_5_n521, po025_driver);
	BUFX2 g_po119 (po119_driver, po119);
	INVX1 g_not_n409 (n409, not_n409);
	INVX1 g_not_n1325_2 (n1325, not_n1325_2);
	AND2X1 g_and_pi079_not_pi136_6 (not_pi136_6, pi079, and_pi079_not_pi136_6);
	AND2X1 g_and_not_n309_not_n335 (not_n309, not_n335, and_not_n309_not_n335);
	BUFX2 g_n448 (and_not_pi016_0_pi054, n448);
	INVX1 g_not_n588 (n588, not_n588);
	INVX1 g_not_n811 (n811, not_n811);
	AND2X1 g_and_not_n850_not_n852 (not_n850, not_n852, and_not_n850_not_n852);
	AND2X1 g_and_pi082_not_n589 (not_n589, pi082, and_pi082_not_n589);
	INVX1 g_not_pi018_2 (pi018, not_pi018_2);
	INVX1 g_not_n793 (n793, not_n793);
	INVX1 g_not_pi138_2 (pi138, not_pi138_2);
	INVX1 g_not_pi129_8235430 (pi129, not_pi129_8235430);
	BUFX2 g_n291 (and_not_pi013_not_pi014, n291);
	INVX1 g_not_n1089 (n1089, not_n1089);
	BUFX2 g_n1209 (and_not_n1205_not_n1208, n1209);
	AND2X1 g_and_not_pi106_5_not_n906 (not_pi106_5, not_n906, and_not_pi106_5_not_n906);
	AND2X1 g_and_pi040_pi082 (pi082, pi040, and_pi040_pi082);
	BUFX2 g_po139_driver (and_pi057_not_pi129_19862745642600749547712274393418170162428858902995921035634302679520490, po139_driver);
	BUFX2 g_po001 (po001_driver, po001);
	BUFX2 g_n1552 (and_pi088_pi138, n1552);
	BUFX2 g_n1252 (and_n1250_n1251, n1252);
	AND2X1 g_and_n445_n463 (n445, n463, and_n445_n463);
	INVX1 g_not_pi111 (pi111, not_pi111);
	AND2X1 g_and_not_pi129_35561530251773635572553173835655155124070416738520070_not_n1405 (not_pi129_35561530251773635572553173835655155124070416738520070, not_n1405, and_not_pi129_35561530251773635572553173835655155124070416738520070_not_n1405);
	AND2X1 g_and_not_pi136_4_not_n1450 (not_pi136_4, not_n1450, and_not_pi136_4_not_n1450);
	INVX1 g_not_pi109_6 (pi109, not_pi109_6);
	BUFX2 g_n827 (and_not_pi129_2326305139872070_not_n826, n827);
	INVX1 g_not_n897 (n897, not_n897);
	BUFX2 g_n451 (and_not_pi005_2_n450, n451);
	INVX1 g_not_n1340 (n1340, not_n1340);
	BUFX2 g_n422 (and_n420_n421, n422);
	BUFX2 g_n1567 (and_not_n1565_not_n1566, n1567);
	INVX1 g_not_pi129_405362155971443868320658661090166738008752222510120837461924544480010 (pi129, not_pi129_405362155971443868320658661090166738008752222510120837461924544480010);
	AND2X1 g_and_not_pi129_6_not_n483 (not_pi129_6, not_n483, and_not_pi129_6_not_n483);
	INVX1 g_not_n989 (n989, not_n989);
	BUFX2 g_n1347 (and_not_pi062_not_pi138_1, n1347);
	BUFX2 g_n1601 (and_n1583_n1600, n1601);
	INVX1 g_not_n741 (n741, not_n741);
	BUFX2 g_n569 (and_n399_n568, n569);
	BUFX2 g_n947 (and_pi082_not_n390, n947);
	AND2X1 g_and_n1251_n1291 (n1251, n1291, and_n1251_n1291);
	INVX1 g_not_pi096_3 (pi096, not_pi096_3);
	INVX1 g_not_pi050_1 (pi050, not_pi050_1);
	AND2X1 g_and_pi031_pi109 (pi031, pi109, and_pi031_pi109);
	BUFX2 g_n366 (and_n312_n357, n366);
	BUFX2 g_n420 (and_n341_n419, n420);
	AND2X1 g_and_not_pi129_168830552257994114252669163302859949191483641195385604940410056010_n1604 (not_pi129_168830552257994114252669163302859949191483641195385604940410056010, n1604, and_not_pi129_168830552257994114252669163302859949191483641195385604940410056010_n1604);
	BUFX2 g_n885 (and_not_n883_not_n884, n885);
	AND2X1 g_and_pi142_n1386 (pi142, n1386, and_pi142_n1386);
	INVX1 g_not_pi024_3 (pi024, not_pi024_3);
	INVX1 g_not_pi097 (pi097, not_pi097);
	AND2X1 g_and_not_pi129_7490483309651862334944941026945644936490_not_n1233 (not_n1233, not_pi129_7490483309651862334944941026945644936490, and_not_pi129_7490483309651862334944941026945644936490_not_n1233);
	BUFX2 g_n421 (and_not_pi021_1_n300, n421);
	AND2X1 g_and_not_pi129_3_not_n437 (not_pi129_3, not_n437, and_not_pi129_3_not_n437);
	AND2X1 g_and_not_pi045_1_n384 (n384, not_pi045_1, and_not_pi045_1_n384);
	BUFX2 g_n592 (and_not_n590_not_n591, n592);
	BUFX2 g_n1348 (and_not_n1346_not_n1347, n1348);
	AND2X1 g_and_not_pi027_3430_n1529 (not_pi027_3430, n1529, and_not_pi027_3430_n1529);
	BUFX2 g_n754 (and_not_pi027_1_not_pi085_3, n754);
	AND2X1 g_and_not_n1399_not_n1400 (not_n1400, not_n1399, and_not_n1399_not_n1400);
	BUFX2 g_n500 (and_pi011_n459, n500);
	BUFX2 g_n1498 (and_not_n1496_not_n1497, n1498);
	BUFX2 g_n349 (and_n344_n348, n349);
	AND2X1 g_and_not_pi040_n390 (n390, not_pi040, and_not_pi040_n390);
	BUFX2 g_n643 (and_not_pi044_0_n401, n643);
	BUFX2 g_po035_driver (and_not_pi129_403536070_not_n660, po035_driver);
	INVX1 g_not_pi129_541169560379521116689596608490 (pi129, not_pi129_541169560379521116689596608490);
	AND2X1 g_and_n301_n302 (n302, n301, and_n301_n302);
	INVX1 g_not_n1164_0 (n1164, not_n1164_0);
	INVX1 g_not_pi043_1 (pi043, not_pi043_1);
	AND2X1 g_and_n754_n787 (n754, n787, and_n754_n787);
	INVX1 g_not_pi014_1 (pi014, not_pi014_1);
	BUFX2 g_n368 (and_not_pi009_0_not_n367, n368);
	AND2X1 g_and_n341_n419 (n341, n419, and_n341_n419);
	BUFX2 g_n674 (and_n448_n673, n674);
	BUFX2 g_n427 (and_not_pi113_n426, n427);
	BUFX2 g_n833 (and_not_n831_not_n832, n833);
	BUFX2 g_n1111 (and_n638_n1110, n1111);
	INVX1 g_not_pi004 (pi004, not_pi004);
	AND2X1 g_and_not_n1515_not_n1516 (not_n1516, not_n1515, and_not_n1515_not_n1516);
	AND2X1 g_and_not_pi129_3788186922656647816827176259430_not_n1060 (not_pi129_3788186922656647816827176259430, not_n1060, and_not_pi129_3788186922656647816827176259430_not_n1060);
	AND2X1 g_and_n550_n551 (n551, n550, and_n550_n551);
	INVX1 g_not_n1007 (n1007, not_n1007);
	AND2X1 g_and_pi034_pi109 (pi034, pi109, and_pi034_pi109);
	INVX1 g_not_n1060 (n1060, not_n1060);
	BUFX2 g_n1083 (and_n379_not_n1082, n1083);
	INVX1 g_not_n1177 (n1177, not_n1177);
	INVX1 g_not_n911 (n911, not_n911);
	BUFX2 g_n1326 (and_pi078_not_n1325, n1326);
	INVX1 g_not_n1438 (n1438, not_n1438);
	AND2X1 g_and_n448_n524 (n524, n448, and_n448_n524);
	INVX1 g_not_pi129_657123623635342801395430 (pi129, not_pi129_657123623635342801395430);
	AND2X1 g_and_not_pi026_5_pi027 (pi027, not_pi026_5, and_not_pi026_5_pi027);
	AND2X1 g_and_not_pi110_1_not_n761 (not_pi110_1, not_n761, and_not_pi110_1_not_n761);
	INVX1 g_not_pi027 (pi027, not_pi027);
	BUFX2 g_n1613 (and_not_pi054_8235430_pi118, n1613);
	BUFX2 g_n388 (and_not_pi038_not_pi050, n388);
	INVX1 g_not_n1503 (n1503, not_n1503);
	BUFX2 g_n377 (and_not_pi129_0_not_n376, n377);
	AND2X1 g_and_n748_n750 (n750, n748, and_n748_n750);
	BUFX2 g_n1124 (and_not_n1119_not_n1123, n1124);
	INVX1 g_not_n1558 (n1558, not_n1558);
	AND2X1 g_and_not_pi136_5_not_n1461 (not_n1461, not_pi136_5, and_not_pi136_5_not_n1461);
	AND2X1 g_and_not_pi129_248930711762415449007872216849586085868492917169640490_not_n1409 (not_pi129_248930711762415449007872216849586085868492917169640490, not_n1409, and_not_pi129_248930711762415449007872216849586085868492917169640490_not_n1409);
	BUFX2 g_n1469 (and_pi138_not_n1468, n1469);
	BUFX2 g_n850 (and_not_pi085_6_not_n849, n850);
	BUFX2 g_n1474 (and_not_pi069_0_pi136, n1474);
	BUFX2 g_n436 (and_pi004_not_pi054, n436);
	BUFX2 g_n688 (and_not_pi047_1_n568, n688);
	INVX1 g_not_n726_1 (n726, not_n726_1);
	BUFX2 g_po132 (po132_driver, po132);
	BUFX2 g_n1507 (and_pi137_not_n1506, n1507);
	AND2X1 g_and_not_n727_not_n728 (not_n728, not_n727, and_not_n727_not_n728);
	AND2X1 g_and_pi017_not_pi054_70 (pi017, not_pi054_70, and_pi017_not_pi054_70);
	BUFX2 g_po092_driver (or_pi129_n1322, po092_driver);
	INVX1 g_not_pi106_8 (pi106, not_pi106_8);
	BUFX2 g_n930 (and_n927_n929, n930);
	BUFX2 g_po063 (po063_driver, po063);
	BUFX2 g_n386 (and_n382_n385, n386);
	INVX1 g_not_n1147 (n1147, not_n1147);
	AND2X1 g_and_pi136_not_n1536 (not_n1536, pi136, and_pi136_not_n1536);
	INVX1 g_not_pi062 (pi062, not_pi062);
	INVX1 g_not_pi106_3 (pi106, not_pi106_3);
	AND2X1 g_and_not_n325_not_n327 (not_n327, not_n325, and_not_n325_not_n327);
	BUFX2 g_n426 (and_pi000_not_pi123, n426);
	INVX1 g_not_pi129_4599865365447399609768010 (pi129, not_pi129_4599865365447399609768010);
	BUFX2 g_n622 (and_n450_n621, n622);
	AND2X1 g_and_not_pi129_541169560379521116689596608490_not_n1044 (not_pi129_541169560379521116689596608490, not_n1044, and_not_pi129_541169560379521116689596608490_not_n1044);
	BUFX2 g_po091_driver (or_pi129_n1318, po091_driver);
	INVX1 g_not_n582 (n582, not_n582);
	AND2X1 g_and_not_n794_not_n795 (not_n795, not_n794, and_not_n794_not_n795);
	INVX1 g_not_n1271 (n1271, not_n1271);
	INVX1 g_not_n1136 (n1136, not_n1136);
	BUFX2 g_n1032 (and_n379_not_n1031, n1032);
	AND2X1 g_and_pi088_pi138 (pi088, pi138, and_pi088_pi138);
	AND2X1 g_and_not_pi046_0_not_pi050_0 (not_pi050_0, not_pi046_0, and_not_pi046_0_not_pi050_0);
	AND2X1 g_and_not_pi024_not_pi049 (not_pi049, not_pi024, and_not_pi024_not_pi049);
	BUFX2 g_n1144 (and_pi058_pi116, n1144);
	BUFX2 g_n363 (and_pi007_n357, n363);
	BUFX2 g_n446 (and_n444_n445, n446);
	AND2X1 g_and_not_n628_not_n634 (not_n628, not_n634, and_not_n628_not_n634);
	BUFX2 g_n796 (and_not_n794_not_n795, n796);
	BUFX2 g_n1173 (and_not_n1168_not_n1172, n1173);
	AND2X1 g_and_not_pi027_70_not_n1198 (not_pi027_70, not_n1198, and_not_pi027_70_not_n1198);
	AND2X1 g_and_not_pi137_10_not_n1560 (not_n1560, not_pi137_10, and_not_pi137_10_not_n1560);
	INVX1 g_not_pi129_85383234134508499009700170379408027452893070589186688070 (pi129, not_pi129_85383234134508499009700170379408027452893070589186688070);
	AND2X1 g_and_not_pi026_24010_not_n1230 (not_n1230, not_pi026_24010, and_not_pi026_24010_not_n1230);
	INVX1 g_not_pi026 (pi026, not_pi026);
	INVX1 g_not_n730 (n730, not_n730);
	INVX1 g_not_n894 (n894, not_n894);
	BUFX2 g_po029_driver (and_not_pi003_9_n566, po029_driver);
	BUFX2 g_n1411 (and_pi082_not_pi137_3, n1411);
	BUFX2 g_n853 (and_not_n850_not_n852, n853);
	INVX1 g_not_n1083 (n1083, not_n1083);
	AND2X1 g_and_not_pi070_0_not_pi138_70 (not_pi070_0, not_pi138_70, and_not_pi070_0_not_pi138_70);
	INVX1 g_not_pi009_1 (pi009, not_pi009_1);
	BUFX2 g_n838 (and_pi029_not_pi116_5, n838);
	AND2X1 g_and_n934_n1131 (n1131, n934, and_n934_n1131);
	AND2X1 g_and_not_pi112_0_not_n1421_1 (not_pi112_0, not_n1421_1, and_not_pi112_0_not_n1421_1);
	BUFX2 g_po077_driver (or_pi129_n1253, po077_driver);
	AND2X1 g_and_not_pi129_16284135979104490_not_n858 (not_pi129_16284135979104490, not_n858, and_not_pi129_16284135979104490_not_n858);
	INVX1 g_not_n1171 (n1171, not_n1171);
	INVX1 g_not_n1523 (n1523, not_n1523);
	INVX1 g_not_n1594 (n1594, not_n1594);
	INVX1 g_not_n906 (n906, not_n906);
	BUFX2 g_po106 (po106_driver, po106);
	BUFX2 g_n1598 (and_not_pi129_24118650322570587750381309043265707027354805885055086420058579430_not_n1597, n1598);
	INVX1 g_not_pi012_0 (pi012, not_pi012_0);
	AND2X1 g_and_not_pi003_138412872010_n1185 (not_pi003_138412872010, n1185, and_not_pi003_138412872010_n1185);
	BUFX2 g_n1377 (and_pi086_not_n1325_5, n1377);
	BUFX2 g_n830 (and_pi097_not_pi110_3, n830);
	INVX1 g_not_pi109_2 (pi109, not_pi109_2);
	AND2X1 g_and_not_pi002_3_n399 (n399, not_pi002_3, and_not_pi002_3_n399);
	AND2X1 g_and_pi082_not_n1101 (pi082, not_n1101, and_pi082_not_n1101);
	BUFX2 g_n1458 (and_pi037_n1360, n1458);
	AND2X1 g_and_pi024_pi082 (pi024, pi082, and_pi024_pi082);
	BUFX2 g_n944 (and_pi039_not_n943, n944);
	INVX1 g_not_pi138_7 (pi138, not_pi138_7);
	AND2X1 g_and_n583_n704 (n704, n583, and_n583_n704);
	BUFX2 g_n695 (and_not_n691_not_n694, n695);
	INVX1 g_not_pi024_2 (pi024, not_pi024_2);
	INVX1 g_not_n842 (n842, not_n842);
	BUFX2 g_n1401 (and_not_n1399_not_n1400, n1401);
	BUFX2 g_n1310 (and_not_n1308_not_n1309, n1310);
	AND2X1 g_and_not_pi051_0_n736 (not_pi051_0, n736, and_not_pi051_0_n736);
	BUFX2 g_n1203 (and_not_pi129_152867006319425761937651857692768264010_not_n1202, n1203);
	BUFX2 g_n520 (and_not_n511_not_n519, n520);
	INVX1 g_not_pi075 (pi075, not_pi075);
	INVX1 g_not_n969 (n969, not_n969);
	BUFX2 g_po075_driver (or_n1237_n1238, po075_driver);
	AND2X1 g_and_not_n764_not_n765 (not_n764, not_n765, and_not_n764_not_n765);
	AND2X1 g_and_not_pi058_5_not_pi110_4 (not_pi058_5, not_pi110_4, and_not_pi058_5_not_pi110_4);
	AND2X1 g_and_not_pi053_5_not_n1148 (not_pi053_5, not_n1148, and_not_pi053_5_not_n1148);
	AND2X1 g_and_pi027_n1182 (n1182, pi027, and_pi027_n1182);
	INVX1 g_not_n1325_0 (n1325, not_n1325_0);
	BUFX2 g_n1367 (and_not_n1365_not_n1366, n1367);
	INVX1 g_not_n1128 (n1128, not_n1128);
	INVX1 g_not_n1327 (n1327, not_n1327);
	AND2X1 g_and_n1412_n1413 (n1412, n1413, and_n1412_n1413);
	AND2X1 g_and_not_pi005_0_not_pi006_1 (not_pi006_1, not_pi005_0, and_not_pi005_0_not_pi006_1);
	BUFX2 g_n1492 (and_not_pi137_6_not_n1491, n1492);
	BUFX2 g_n692 (and_n584_n650, n692);
	AND2X1 g_and_not_pi106_0_not_n871 (not_n871, not_pi106_0, and_not_pi106_0_not_n871);
	INVX1 g_not_n1247_3 (n1247, not_n1247_3);
	AND2X1 g_and_n448_n451 (n451, n448, and_n448_n451);
	BUFX2 g_n403 (and_not_pi038_0_not_pi040_0, n403);
	INVX1 g_not_pi054_7 (pi054, not_pi054_7);
	INVX1 g_not_n924 (n924, not_n924);
	INVX1 g_not_pi054_168070 (pi054, not_pi054_168070);
	BUFX2 g_n869 (and_pi030_pi109, n869);
	AND2X1 g_and_n705_n1106 (n1106, n705, and_n705_n1106);
	AND2X1 g_and_n331_n332 (n332, n331, and_n331_n332);
	INVX1 g_not_pi085_5 (pi085, not_pi085_5);
	BUFX2 g_n1541 (and_not_pi136_24010_not_n1540, n1541);
	AND2X1 g_and_n638_n639 (n638, n639, and_n638_n639);
	BUFX2 g_n1420 (and_not_pi110_6_n1419, n1420);
	BUFX2 g_n1545 (and_pi081_not_pi138_1176490, n1545);
	AND2X1 g_and_n448_n673 (n673, n448, and_n448_n673);
	BUFX2 g_n943 (and_pi109_n722, n943);
	INVX1 g_not_n901 (n901, not_n901);
	AND2X1 g_and_not_n910_not_n914 (not_n910, not_n914, and_not_n910_not_n914);
	INVX1 g_not_n751 (n751, not_n751);
	BUFX2 g_n1107 (and_n705_n1106, n1107);
	INVX1 g_not_n761_0 (n761, not_n761_0);
	AND2X1 g_and_not_pi018_0_n449 (n449, not_pi018_0, and_not_pi018_0_n449);
	BUFX2 g_n470 (and_not_pi129_5_not_n469, n470);
	BUFX2 g_n1449 (and_not_pi077_not_pi138_5, n1449);
	AND2X1 g_and_not_pi016_2_n351 (not_pi016_2, n351, and_not_pi016_2_n351);
	INVX1 g_not_pi137 (pi137, not_pi137);
	INVX1 g_not_n1421_1 (n1421, not_n1421_1);
	AND2X1 g_and_not_n782_not_n783 (not_n783, not_n782, and_not_n782_not_n783);
	AND2X1 g_and_pi012_not_pi054_7 (pi012, not_pi054_7, and_pi012_not_pi054_7);
	BUFX2 g_n896 (and_pi092_pi106, n896);
	INVX1 g_not_n810 (n810, not_n810);
	BUFX2 g_n821 (and_n819_n820, n821);
	AND2X1 g_and_not_pi011_2_pi021 (not_pi011_2, pi021, and_not_pi011_2_pi021);
	BUFX2 g_n348 (and_not_pi014_1_n347, n348);
	AND2X1 g_and_pi011_n459 (n459, pi011, and_pi011_n459);
	BUFX2 g_n1034 (and_not_pi045_4_not_n1033, n1034);
	AND2X1 g_and_not_n1164_not_n1166 (not_n1166, not_n1164, and_not_n1164_not_n1166);
	INVX1 g_not_n1220 (n1220, not_n1220);
	BUFX2 g_n1373 (and_not_pi129_43181145673964365640352930977077280875522488490_not_n1372, n1373);
	AND2X1 g_and_n300_n303 (n303, n300, and_n300_n303);
	AND2X1 g_and_not_pi027_2_not_pi053_1 (not_pi053_1, not_pi027_2, and_not_pi027_2_not_pi053_1);
	AND2X1 g_and_n838_n856 (n838, n856, and_n838_n856);
	AND2X1 g_and_not_pi116_6_n843 (not_pi116_6, n843, and_not_pi116_6_n843);
	AND2X1 g_and_n1175_n1182 (n1182, n1175, and_n1175_n1182);
	INVX1 g_not_pi003_57648010 (pi003, not_pi003_57648010);
	BUFX2 g_n702 (and_not_n379_2_not_n701, n702);
	AND2X1 g_and_not_n604_not_n616 (not_n604, not_n616, and_not_n604_not_n616);
	AND2X1 g_and_n291_n344 (n344, n291, and_n291_n344);
	BUFX2 g_n703 (and_pi063_n702, n703);
	INVX1 g_not_pi053_2 (pi053, not_pi053_2);
	INVX1 g_not_pi005_3 (pi005, not_pi005_3);
	BUFX2 g_n1417 (and_not_n1415_not_n1416, n1417);
	INVX1 g_not_pi136_5 (pi136, not_pi136_5);
	BUFX2 g_n568 (and_not_pi041_1_not_pi043_1, n568);
	BUFX2 g_n651 (and_n390_n650, n651);
	BUFX2 g_n341 (and_not_pi011_0_not_pi012_1, n341);
	INVX1 g_not_pi116_2 (pi116, not_pi116_2);
	BUFX2 g_n338 (and_not_n307_not_n337, n338);
	INVX1 g_not_n1519 (n1519, not_n1519);
	INVX1 g_not_pi058_9 (pi058, not_pi058_9);
	AND2X1 g_and_pi009_n369 (n369, pi009, and_pi009_n369);
	BUFX2 g_po115 (po115_driver, po115);
	BUFX2 g_n1362 (and_not_n1359_not_n1361, n1362);
	AND2X1 g_and_pi098_not_n1386_5 (not_n1386_5, pi098, and_pi098_not_n1386_5);
	AND2X1 g_and_not_pi140_n1249 (n1249, not_pi140, and_not_pi140_n1249);
	BUFX2 g_n615 (and_n611_n614, n615);
	INVX1 g_not_pi017 (pi017, not_pi017);
	BUFX2 g_n1199 (and_not_pi027_70_not_n1198, n1199);
	BUFX2 g_n1251 (and_not_pi138_0_n1246, n1251);
	BUFX2 g_n868 (and_pi089_pi106, n868);
	INVX1 g_not_n310 (n310, not_n310);
	INVX1 g_not_pi027_8 (pi027, not_pi027_8);
	INVX1 g_not_pi109_7 (pi109, not_pi109_7);
	BUFX2 g_n1520 (and_not_pi137_8_not_n1519, n1520);
	BUFX2 g_n779 (and_n776_n778, n779);
	BUFX2 g_n1382 (and_pi140_n1325, n1382);
	INVX1 g_not_n368 (n368, not_n368);
	BUFX2 g_n616 (and_n609_n615, n616);
	AND2X1 g_and_pi109_n722 (n722, pi109, and_pi109_n722);
	INVX1 g_not_n967 (n967, not_n967);
	INVX1 g_not_n1304 (n1304, not_n1304);
	BUFX2 g_n1486 (and_pi033_pi136, n1486);
	AND2X1 g_and_n385_n1035 (n1035, n385, and_n385_n1035);
	INVX1 g_not_n1115 (n1115, not_n1115);
	OR2X1 g_or_n1520_n1527 (n1527, n1520, or_n1520_n1527);
	AND2X1 g_and_not_n717_not_n719 (not_n719, not_n717, and_not_n717_not_n719);
	INVX1 g_not_pi136_2 (pi136, not_pi136_2);
	INVX1 g_not_pi016_0 (pi016, not_pi016_0);
	INVX1 g_not_pi011 (pi011, not_pi011);
	INVX1 g_not_n681 (n681, not_n681);
	INVX1 g_not_pi112_0 (pi112, not_pi112_0);
	AND2X1 g_and_not_n423_n424 (n424, not_n423, and_not_n423_n424);
	INVX1 g_not_n379_490 (n379, not_n379_490);
	BUFX2 g_po019 (po019_driver, po019);
	BUFX2 g_n458 (and_pi006_not_pi054_1, n458);
	INVX1 g_not_pi129_6782230728490 (pi129, not_pi129_6782230728490);
	BUFX2 g_n1061 (and_not_pi129_3788186922656647816827176259430_not_n1060, n1061);
	INVX1 g_not_n1353 (n1353, not_n1353);
	AND2X1 g_and_not_pi007_10_not_pi009_6 (not_pi009_6, not_pi007_10, and_not_pi007_10_not_pi009_6);
	BUFX2 g_po074_driver (and_not_pi003_47475615099430_n1234, po074_driver);
	INVX1 g_not_pi020_0 (pi020, not_pi020_0);
	BUFX2 g_n841 (and_not_n836_not_n840, n841);
	BUFX2 g_n724 (and_not_pi095_not_pi100, n724);
	AND2X1 g_and_not_pi047_2_n407 (n407, not_pi047_2, and_not_pi047_2_n407);
	INVX1 g_not_n1180 (n1180, not_n1180);
	INVX1 g_not_n590 (n590, not_n590);
	AND2X1 g_and_not_n1504_not_n1505 (not_n1504, not_n1505, and_not_n1504_not_n1505);
	BUFX2 g_n316 (and_not_n314_not_n315, n316);
	INVX1 g_not_pi138 (pi138, not_pi138);
	BUFX2 g_n477 (and_n448_n476, n477);
	INVX1 g_not_n693 (n693, not_n693);
	AND2X1 g_and_not_pi026_2_n713 (n713, not_pi026_2, and_not_pi026_2_n713);
	BUFX2 g_n1153 (and_not_pi129_3119734822845423713013303218219760490_not_n1152, n1153);
	INVX1 g_not_pi015_2 (pi015, not_pi015_2);
	BUFX2 g_po084_driver (or_pi129_n1288, po084_driver);
	BUFX2 g_n1151 (and_not_pi116_6_n843, n1151);
	BUFX2 g_n1128 (and_pi082_not_n1127, n1128);
	AND2X1 g_and_pi027_not_n739 (not_n739, pi027, and_pi027_not_n739);
	INVX1 g_not_pi137_0 (pi137, not_pi137_0);
	BUFX2 g_n488 (and_not_pi017_4_not_pi018_2, n488);
	INVX1 g_not_pi136_1176490 (pi136, not_pi136_1176490);
	AND2X1 g_and_not_pi023_pi055 (not_pi023, pi055, and_not_pi023_pi055);
	INVX1 g_not_n1396 (n1396, not_n1396);
	AND2X1 g_and_pi099_pi106 (pi106, pi099, and_pi099_pi106);
	AND2X1 g_and_pi082_not_n1069 (pi082, not_n1069, and_pi082_not_n1069);
	AND2X1 g_and_pi098_pi138 (pi138, pi098, and_pi098_pi138);
	INVX1 g_not_pi109_5 (pi109, not_pi109_5);
	BUFX2 g_n995 (and_pi072_n994, n995);
	AND2X1 g_and_not_pi136_not_pi137_1 (not_pi136, not_pi137_1, and_not_pi136_not_pi137_1);
	AND2X1 g_and_n1244_n1246 (n1246, n1244, and_n1244_n1246);
	INVX1 g_not_n1481 (n1481, not_n1481);
	INVX1 g_not_n1554 (n1554, not_n1554);
	AND2X1 g_and_pi054_not_n1595 (not_n1595, pi054, and_pi054_not_n1595);
	AND2X1 g_and_n388_n390 (n388, n390, and_n388_n390);
	INVX1 g_not_n735 (n735, not_n735);
	INVX1 g_not_n1521 (n1521, not_n1521);
	BUFX2 g_n295 (and_not_pi008_n294, n295);
	AND2X1 g_and_n343_n349 (n349, n343, and_n343_n349);
	BUFX2 g_po078_driver (or_pi129_n1258, po078_driver);
	BUFX2 g_n1286 (and_not_pi143_0_n1249, n1286);
	BUFX2 g_n1481 (and_pi090_n1249, n1481);
	INVX1 g_not_n1056 (n1056, not_n1056);
	BUFX2 g_n1125 (and_not_pi050_4_not_n1124, n1125);
	AND2X1 g_and_not_n1308_not_n1309 (not_n1309, not_n1308, and_not_n1308_not_n1309);
	BUFX2 g_n337 (and_pi054_not_n336, n337);
	BUFX2 g_n856 (and_pi026_n855, n856);
	BUFX2 g_n963 (and_not_n959_n962, n963);
	INVX1 g_not_n738 (n738, not_n738);
	AND2X1 g_and_not_pi041_1_not_pi043_1 (not_pi041_1, not_pi043_1, and_not_pi041_1_not_pi043_1);
	INVX1 g_not_pi007_7 (pi007, not_pi007_7);
	AND2X1 g_and_n743_n755 (n743, n755, and_n743_n755);
	AND2X1 g_and_not_n831_not_n832 (not_n832, not_n831, and_not_n831_not_n832);
	INVX1 g_not_n1164 (n1164, not_n1164);
	INVX1 g_not_pi118 (pi118, not_pi118);
	INVX1 g_not_n912 (n912, not_n912);
	INVX1 g_not_n309 (n309, not_n309);
	BUFX2 g_n1060 (and_n1054_n1059, n1060);
	AND2X1 g_and_not_n889_not_n893 (not_n893, not_n889, and_not_n889_not_n893);
	AND2X1 g_and_not_n435_not_n436 (not_n436, not_n435, and_not_n435_not_n436);
	BUFX2 g_n1472 (and_not_n1470_not_n1471, n1472);
	AND2X1 g_and_pi094_n1324 (pi094, n1324, and_pi094_n1324);
	BUFX2 g_n414 (and_not_n397_not_n413, n414);
	INVX1 g_not_n726 (n726, not_n726);
	INVX1 g_not_n724 (n724, not_n724);
	AND2X1 g_and_not_n440_not_n454 (not_n440, not_n454, and_not_n440_not_n454);
	AND2X1 g_and_pi116_n1165 (pi116, n1165, and_pi116_n1165);
	BUFX2 g_n1297 (and_n1251_n1296, n1297);
	BUFX2 g_n506 (and_n503_n505, n506);
	INVX1 g_not_pi137_6 (pi137, not_pi137_6);
	AND2X1 g_and_pi009_not_pi054_4 (not_pi054_4, pi009, and_pi009_not_pi054_4);
	INVX1 g_not_n803 (n803, not_n803);
	INVX1 g_not_n727 (n727, not_n727);
	AND2X1 g_and_pi123_n1236 (n1236, pi123, and_pi123_n1236);
	INVX1 g_not_pi003_3430 (pi003, not_pi003_3430);
	BUFX2 g_n532 (and_not_pi129_10_not_n531, n532);
	BUFX2 g_po020_driver (and_not_pi003_0_n456, po020_driver);
	BUFX2 g_n664 (and_not_pi021_3_pi054, n664);
	BUFX2 g_n546 (and_n448_n545, n546);

endmodule
