module adder(
    N1,
    N2,
    N3,
    N4,
    N5,
    N6,
    N7,
    N8,
    N9,
    N10,
    N11,
    N12,
    N13,
    N14,
    N15,
    N16,
    N17,
    N18,
    N19,
    N20,
    N21,
    N22,
    N23,
    N24,
    N25,
    N26,
    N27,
    N28,
    N29,
    N30,
    N31,
    N32,
    N33,
    N34,
    N35,
    N36,
    N37,
    N38,
    N39,
    N40,
    N41,
    N42,
    N43,
    N44,
    N45,
    N46,
    N47,
    N48,
    N49,
    N50,
    N51,
    N52,
    N53,
    N54,
    N55,
    N56,
    N57,
    N58,
    N59,
    N60,
    N61,
    N62,
    N63,
    N64,
    N65,
    N66,
    N67,
    N68,
    N69,
    N70,
    N71,
    N72,
    N73,
    N74,
    N75,
    N76,
    N77,
    N78,
    N79,
    N80,
    N81,
    N82,
    N83,
    N84,
    N85,
    N86,
    N87,
    N88,
    N89,
    N90,
    N91,
    N92,
    N93,
    N94,
    N95,
    N96,
    N97,
    N98,
    N99,
    N100,
    N101,
    N102,
    N103,
    N104,
    N105,
    N106,
    N107,
    N108,
    N109,
    N110,
    N111,
    N112,
    N113,
    N114,
    N115,
    N116,
    N117,
    N118,
    N119,
    N120,
    N121,
    N122,
    N123,
    N124,
    N125,
    N126,
    N127,
    N128,
    N129,
    N130,
    N131,
    N132,
    N133,
    N134,
    N135,
    N136,
    N137,
    N138,
    N139,
    N140,
    N141,
    N142,
    N143,
    N144,
    N145,
    N146,
    N147,
    N148,
    N149,
    N150,
    N151,
    N152,
    N153,
    N154,
    N155,
    N156,
    N157,
    N158,
    N159,
    N160,
    N161,
    N162,
    N163,
    N164,
    N165,
    N166,
    N167,
    N168,
    N169,
    N170,
    N171,
    N172,
    N173,
    N174,
    N175,
    N176,
    N177,
    N178,
    N179,
    N180,
    N181,
    N182,
    N183,
    N184,
    N185,
    N186,
    N187,
    N188,
    N189,
    N190,
    N191,
    N192,
    N193,
    N194,
    N195,
    N196,
    N197,
    N198,
    N199,
    N200,
    N201,
    N202,
    N203,
    N204,
    N205,
    N206,
    N207,
    N208,
    N209,
    N210,
    N211,
    N212,
    N213,
    N214,
    N215,
    N216,
    N217,
    N218,
    N219,
    N220,
    N221,
    N222,
    N223,
    N224,
    N225,
    N226,
    N227,
    N228,
    N229,
    N230,
    N231,
    N232,
    N233,
    N234,
    N235,
    N236,
    N237,
    N238,
    N239,
    N240,
    N241,
    N242,
    N243,
    N244,
    N245,
    N246,
    N247,
    N248,
    N249,
    N250,
    N251,
    N252,
    N253,
    N254,
    N255,
    N256,
    N257,
    N258,
    N259,
    N260,
    N261,
    N262,
    N263,
    N264,
    N265,
    N266,
    N267,
    N268,
    N269,
    N270,
    N271,
    N272,
    N273,
    N274,
    N275,
    N276,
    N277,
    N278,
    N279,
    N280,
    N281,
    N282,
    N283,
    N284,
    N285,
    N286,
    N287,
    N288,
    N289,
    N290,
    N291,
    N292,
    N293,
    N294,
    N295,
    N296,
    N297,
    N298,
    N299,
    N300,
    N301,
    N302,
    N303,
    N304,
    N305,
    N306,
    N307,
    N308,
    N309,
    N310,
    N311,
    N312,
    N313,
    N314,
    N315,
    N316,
    N317,
    N318,
    N319,
    N320,
    N321,
    N322,
    N323,
    N324,
    N325,
    N326,
    N327,
    N328,
    N329,
    N330,
    N331,
    N332,
    N333,
    N334,
    N335,
    N336,
    N337,
    N338,
    N339,
    N340,
    N341,
    N342,
    N343,
    N344,
    N345,
    N346,
    N347,
    N348,
    N349,
    N350,
    N351,
    N352,
    N353,
    N354,
    N355,
    N356,
    N357,
    N358,
    N359,
    N360,
    N361,
    N362,
    N363,
    N364,
    N365,
    N366,
    N367,
    N368,
    N369,
    N370,
    N371,
    N372,
    N373,
    N374,
    N375,
    N376,
    N377,
    N378,
    N379,
    N380,
    N381,
    N382,
    N383,
    N384,
    N385);
    input N1;
    input N2;
    input N3;
    input N4;
    input N5;
    input N6;
    input N7;
    input N8;
    input N9;
    input N10;
    input N11;
    input N12;
    input N13;
    input N14;
    input N15;
    input N16;
    input N17;
    input N18;
    input N19;
    input N20;
    input N21;
    input N22;
    input N23;
    input N24;
    input N25;
    input N26;
    input N27;
    input N28;
    input N29;
    input N30;
    input N31;
    input N32;
    input N33;
    input N34;
    input N35;
    input N36;
    input N37;
    input N38;
    input N39;
    input N40;
    input N41;
    input N42;
    input N43;
    input N44;
    input N45;
    input N46;
    input N47;
    input N48;
    input N49;
    input N50;
    input N51;
    input N52;
    input N53;
    input N54;
    input N55;
    input N56;
    input N57;
    input N58;
    input N59;
    input N60;
    input N61;
    input N62;
    input N63;
    input N64;
    input N65;
    input N66;
    input N67;
    input N68;
    input N69;
    input N70;
    input N71;
    input N72;
    input N73;
    input N74;
    input N75;
    input N76;
    input N77;
    input N78;
    input N79;
    input N80;
    input N81;
    input N82;
    input N83;
    input N84;
    input N85;
    input N86;
    input N87;
    input N88;
    input N89;
    input N90;
    input N91;
    input N92;
    input N93;
    input N94;
    input N95;
    input N96;
    input N97;
    input N98;
    input N99;
    input N100;
    input N101;
    input N102;
    input N103;
    input N104;
    input N105;
    input N106;
    input N107;
    input N108;
    input N109;
    input N110;
    input N111;
    input N112;
    input N113;
    input N114;
    input N115;
    input N116;
    input N117;
    input N118;
    input N119;
    input N120;
    input N121;
    input N122;
    input N123;
    input N124;
    input N125;
    input N126;
    input N127;
    input N128;
    input N129;
    input N130;
    input N131;
    input N132;
    input N133;
    input N134;
    input N135;
    input N136;
    input N137;
    input N138;
    input N139;
    input N140;
    input N141;
    input N142;
    input N143;
    input N144;
    input N145;
    input N146;
    input N147;
    input N148;
    input N149;
    input N150;
    input N151;
    input N152;
    input N153;
    input N154;
    input N155;
    input N156;
    input N157;
    input N158;
    input N159;
    input N160;
    input N161;
    input N162;
    input N163;
    input N164;
    input N165;
    input N166;
    input N167;
    input N168;
    input N169;
    input N170;
    input N171;
    input N172;
    input N173;
    input N174;
    input N175;
    input N176;
    input N177;
    input N178;
    input N179;
    input N180;
    input N181;
    input N182;
    input N183;
    input N184;
    input N185;
    input N186;
    input N187;
    input N188;
    input N189;
    input N190;
    input N191;
    input N192;
    input N193;
    input N194;
    input N195;
    input N196;
    input N197;
    input N198;
    input N199;
    input N200;
    input N201;
    input N202;
    input N203;
    input N204;
    input N205;
    input N206;
    input N207;
    input N208;
    input N209;
    input N210;
    input N211;
    input N212;
    input N213;
    input N214;
    input N215;
    input N216;
    input N217;
    input N218;
    input N219;
    input N220;
    input N221;
    input N222;
    input N223;
    input N224;
    input N225;
    input N226;
    input N227;
    input N228;
    input N229;
    input N230;
    input N231;
    input N232;
    input N233;
    input N234;
    input N235;
    input N236;
    input N237;
    input N238;
    input N239;
    input N240;
    input N241;
    input N242;
    input N243;
    input N244;
    input N245;
    input N246;
    input N247;
    input N248;
    input N249;
    input N250;
    input N251;
    input N252;
    input N253;
    input N254;
    input N255;
    input N256;
    output N257;
    output N258;
    output N259;
    output N260;
    output N261;
    output N262;
    output N263;
    output N264;
    output N265;
    output N266;
    output N267;
    output N268;
    output N269;
    output N270;
    output N271;
    output N272;
    output N273;
    output N274;
    output N275;
    output N276;
    output N277;
    output N278;
    output N279;
    output N280;
    output N281;
    output N282;
    output N283;
    output N284;
    output N285;
    output N286;
    output N287;
    output N288;
    output N289;
    output N290;
    output N291;
    output N292;
    output N293;
    output N294;
    output N295;
    output N296;
    output N297;
    output N298;
    output N299;
    output N300;
    output N301;
    output N302;
    output N303;
    output N304;
    output N305;
    output N306;
    output N307;
    output N308;
    output N309;
    output N310;
    output N311;
    output N312;
    output N313;
    output N314;
    output N315;
    output N316;
    output N317;
    output N318;
    output N319;
    output N320;
    output N321;
    output N322;
    output N323;
    output N324;
    output N325;
    output N326;
    output N327;
    output N328;
    output N329;
    output N330;
    output N331;
    output N332;
    output N333;
    output N334;
    output N335;
    output N336;
    output N337;
    output N338;
    output N339;
    output N340;
    output N341;
    output N342;
    output N343;
    output N344;
    output N345;
    output N346;
    output N347;
    output N348;
    output N349;
    output N350;
    output N351;
    output N352;
    output N353;
    output N354;
    output N355;
    output N356;
    output N357;
    output N358;
    output N359;
    output N360;
    output N361;
    output N362;
    output N363;
    output N364;
    output N365;
    output N366;
    output N367;
    output N368;
    output N369;
    output N370;
    output N371;
    output N372;
    output N373;
    output N374;
    output N375;
    output N376;
    output N377;
    output N378;
    output N379;
    output N380;
    output N381;
    output N382;
    output N383;
    output N384;
    output N385;

    // Internal wires
    wire N386;
    wire N387;
    wire N388;
    wire N389;
    wire N390;
    wire N391;
    wire N392;
    wire N393;
    wire N394;
    wire N395;
    wire N396;
    wire N397;
    wire N398;
    wire N399;
    wire N400;
    wire N401;
    wire N402;
    wire N403;
    wire N404;
    wire N405;
    wire N406;
    wire N407;
    wire N408;
    wire N409;
    wire N410;
    wire N411;
    wire N412;
    wire N413;
    wire N414;
    wire N415;
    wire N416;
    wire N417;
    wire N418;
    wire N419;
    wire N420;
    wire N421;
    wire N422;
    wire N423;
    wire N424;
    wire N425;
    wire N426;
    wire N427;
    wire N428;
    wire N429;
    wire N430;
    wire N431;
    wire N432;
    wire N433;
    wire N434;
    wire N435;
    wire N436;
    wire N437;
    wire N438;
    wire N439;
    wire N440;
    wire N441;
    wire N442;
    wire N443;
    wire N444;
    wire N445;
    wire N446;
    wire N447;
    wire N448;
    wire N449;
    wire N450;
    wire N451;
    wire N452;
    wire N453;
    wire N454;
    wire N455;
    wire N456;
    wire N457;
    wire N458;
    wire N459;
    wire N460;
    wire N461;
    wire N462;
    wire N463;
    wire N464;
    wire N465;
    wire N466;
    wire N467;
    wire N468;
    wire N469;
    wire N470;
    wire N471;
    wire N472;
    wire N473;
    wire N474;
    wire N475;
    wire N476;
    wire N477;
    wire N478;
    wire N479;
    wire N480;
    wire N481;
    wire N482;
    wire N483;
    wire N484;
    wire N485;
    wire N486;
    wire N487;
    wire N488;
    wire N489;
    wire N490;
    wire N491;
    wire N492;
    wire N493;
    wire N494;
    wire N495;
    wire N496;
    wire N497;
    wire N498;
    wire N499;
    wire N500;
    wire N501;
    wire N502;
    wire N503;
    wire N504;
    wire N505;
    wire N506;
    wire N507;
    wire N508;
    wire N509;
    wire N510;
    wire N511;
    wire N512;
    wire N513;
    wire N514;
    wire N515;
    wire N516;
    wire N517;
    wire N518;
    wire N519;
    wire N520;
    wire N521;
    wire N522;
    wire N523;
    wire N524;
    wire N525;
    wire N526;
    wire N527;
    wire N528;
    wire N529;
    wire N530;
    wire N531;
    wire N532;
    wire N533;
    wire N534;
    wire N535;
    wire N536;
    wire N537;
    wire N538;
    wire N539;
    wire N540;
    wire N541;
    wire N542;
    wire N543;
    wire N544;
    wire N545;
    wire N546;
    wire N547;
    wire N548;
    wire N549;
    wire N550;
    wire N551;
    wire N552;
    wire N553;
    wire N554;
    wire N555;
    wire N556;
    wire N557;
    wire N558;
    wire N559;
    wire N560;
    wire N561;
    wire N562;
    wire N563;
    wire N564;
    wire N565;
    wire N566;
    wire N567;
    wire N568;
    wire N569;
    wire N570;
    wire N571;
    wire N572;
    wire N573;
    wire N574;
    wire N575;
    wire N576;
    wire N577;
    wire N578;
    wire N579;
    wire N580;
    wire N581;
    wire N582;
    wire N583;
    wire N584;
    wire N585;
    wire N586;
    wire N587;
    wire N588;
    wire N589;
    wire N590;
    wire N591;
    wire N592;
    wire N593;
    wire N594;
    wire N595;
    wire N596;
    wire N597;
    wire N598;
    wire N599;
    wire N600;
    wire N601;
    wire N602;
    wire N603;
    wire N604;
    wire N605;
    wire N606;
    wire N607;
    wire N608;
    wire N609;
    wire N610;
    wire N611;
    wire N612;
    wire N613;
    wire N614;
    wire N615;
    wire N616;
    wire N617;
    wire N618;
    wire N619;
    wire N620;
    wire N621;
    wire N622;
    wire N623;
    wire N624;
    wire N625;
    wire N626;
    wire N627;
    wire N628;
    wire N629;
    wire N630;
    wire N631;
    wire N632;
    wire N633;
    wire N634;
    wire N635;
    wire N636;
    wire N637;
    wire N638;
    wire N639;
    wire N640;
    wire N641;
    wire N642;
    wire N643;
    wire N644;
    wire N645;
    wire N646;
    wire N647;
    wire N648;
    wire N649;
    wire N650;
    wire N651;
    wire N652;
    wire N653;
    wire N654;
    wire N655;
    wire N656;
    wire N657;
    wire N658;
    wire N659;
    wire N660;
    wire N661;
    wire N662;
    wire N663;
    wire N664;
    wire N665;
    wire N666;
    wire N667;
    wire N668;
    wire N669;
    wire N670;
    wire N671;
    wire N672;
    wire N673;
    wire N674;
    wire N675;
    wire N676;
    wire N677;
    wire N678;
    wire N679;
    wire N680;
    wire N681;
    wire N682;
    wire N683;
    wire N684;
    wire N685;
    wire N686;
    wire N687;
    wire N688;
    wire N689;
    wire N690;
    wire N691;
    wire N692;
    wire N693;
    wire N694;
    wire N695;
    wire N696;
    wire N697;
    wire N698;
    wire N699;
    wire N700;
    wire N701;
    wire N702;
    wire N703;
    wire N704;
    wire N705;
    wire N706;
    wire N707;
    wire N708;
    wire N709;
    wire N710;
    wire N711;
    wire N712;
    wire N713;
    wire N714;
    wire N715;
    wire N716;
    wire N717;
    wire N718;
    wire N719;
    wire N720;
    wire N721;
    wire N722;
    wire N723;
    wire N724;
    wire N725;
    wire N726;
    wire N727;
    wire N728;
    wire N729;
    wire N730;
    wire N731;
    wire N732;
    wire N733;
    wire N734;
    wire N735;
    wire N736;
    wire N737;
    wire N738;
    wire N739;
    wire N740;
    wire N741;
    wire N742;
    wire N743;
    wire N744;
    wire N745;
    wire N746;
    wire N747;
    wire N748;
    wire N749;
    wire N750;
    wire N751;
    wire N752;
    wire N753;
    wire N754;
    wire N755;
    wire N756;
    wire N757;
    wire N758;
    wire N759;
    wire N760;
    wire N761;
    wire N762;
    wire N763;
    wire N764;
    wire N765;
    wire N766;
    wire N767;
    wire N768;
    wire N769;
    wire N770;
    wire N771;
    wire N772;
    wire N773;
    wire N774;
    wire N775;
    wire N776;
    wire N777;
    wire N778;
    wire N779;
    wire N780;
    wire N781;
    wire N782;
    wire N783;
    wire N784;
    wire N785;
    wire N786;
    wire N787;
    wire N788;
    wire N789;
    wire N790;
    wire N791;
    wire N792;
    wire N793;
    wire N794;
    wire N795;
    wire N796;
    wire N797;
    wire N798;
    wire N799;
    wire N800;
    wire N801;
    wire N802;
    wire N803;
    wire N804;
    wire N805;
    wire N806;
    wire N807;
    wire N808;
    wire N809;
    wire N810;
    wire N811;
    wire N812;
    wire N813;
    wire N814;
    wire N815;
    wire N816;
    wire N817;
    wire N818;
    wire N819;
    wire N820;
    wire N821;
    wire N822;
    wire N823;
    wire N824;
    wire N825;
    wire N826;
    wire N827;
    wire N828;
    wire N829;
    wire N830;
    wire N831;
    wire N832;
    wire N833;
    wire N834;
    wire N835;
    wire N836;
    wire N837;
    wire N838;
    wire N839;
    wire N840;
    wire N841;
    wire N842;
    wire N843;
    wire N844;
    wire N845;
    wire N846;
    wire N847;
    wire N848;
    wire N849;
    wire N850;
    wire N851;
    wire N852;
    wire N853;
    wire N854;
    wire N855;
    wire N856;
    wire N857;
    wire N858;
    wire N859;
    wire N860;
    wire N861;
    wire N862;
    wire N863;
    wire N864;
    wire N865;
    wire N866;
    wire N867;
    wire N868;
    wire N869;
    wire N870;
    wire N871;
    wire N872;
    wire N873;
    wire N874;
    wire N875;
    wire N876;
    wire N877;
    wire N878;
    wire N879;
    wire N880;
    wire N881;
    wire N882;
    wire N883;
    wire N884;
    wire N885;
    wire N886;
    wire N887;
    wire N888;
    wire N889;
    wire N890;
    wire N891;
    wire N892;
    wire N893;
    wire N894;
    wire N895;
    wire N896;
    wire N897;
    wire N898;
    wire N899;
    wire N900;
    wire N901;
    wire N902;
    wire N903;
    wire N904;
    wire N905;
    wire N906;
    wire N907;
    wire N908;
    wire N909;
    wire N910;
    wire N911;
    wire N912;
    wire N913;
    wire N914;
    wire N915;
    wire N916;
    wire N917;
    wire N918;
    wire N919;
    wire N920;
    wire N921;
    wire N922;
    wire N923;
    wire N924;
    wire N925;
    wire N926;
    wire N927;
    wire N928;
    wire N929;
    wire N930;
    wire N931;
    wire N932;
    wire N933;
    wire N934;
    wire N935;
    wire N936;
    wire N937;
    wire N938;
    wire N939;
    wire N940;
    wire N941;
    wire N942;
    wire N943;
    wire N944;
    wire N945;
    wire N946;
    wire N947;
    wire N948;
    wire N949;
    wire N950;
    wire N951;
    wire N952;
    wire N953;
    wire N954;
    wire N955;
    wire N956;
    wire N957;
    wire N958;
    wire N959;
    wire N960;
    wire N961;
    wire N962;
    wire N963;
    wire N964;
    wire N965;
    wire N966;
    wire N967;
    wire N968;
    wire N969;
    wire N970;
    wire N971;
    wire N972;
    wire N973;
    wire N974;
    wire N975;
    wire N976;
    wire N977;
    wire N978;
    wire N979;
    wire N980;
    wire N981;
    wire N982;
    wire N983;
    wire N984;
    wire N985;
    wire N986;
    wire N987;
    wire N988;
    wire N989;
    wire N990;
    wire N991;
    wire N992;
    wire N993;
    wire N994;
    wire N995;
    wire N996;
    wire N997;
    wire N998;
    wire N999;
    wire N1000;
    wire N1001;
    wire N1002;
    wire N1003;
    wire N1004;
    wire N1005;
    wire N1006;
    wire N1007;
    wire N1008;
    wire N1009;
    wire N1010;
    wire N1011;
    wire N1012;
    wire N1013;
    wire N1014;
    wire N1015;
    wire N1016;
    wire N1017;
    wire N1018;
    wire N1019;
    wire N1020;
    wire N1021;
    wire N1022;
    wire N1023;
    wire N1024;
    wire N1025;
    wire N1026;
    wire N1027;
    wire N1028;
    wire N1029;
    wire N1030;
    wire N1031;
    wire N1032;
    wire N1033;
    wire N1034;
    wire N1035;
    wire N1036;
    wire N1037;
    wire N1038;
    wire N1039;
    wire N1040;
    wire N1041;
    wire N1042;
    wire N1043;
    wire N1044;
    wire N1045;
    wire N1046;
    wire N1047;
    wire N1048;
    wire N1049;
    wire N1050;
    wire N1051;
    wire N1052;
    wire N1053;
    wire N1054;
    wire N1055;
    wire N1056;
    wire N1057;
    wire N1058;
    wire N1059;
    wire N1060;
    wire N1061;
    wire N1062;
    wire N1063;
    wire N1064;
    wire N1065;
    wire N1066;
    wire N1067;
    wire N1068;
    wire N1069;
    wire N1070;
    wire N1071;
    wire N1072;
    wire N1073;
    wire N1074;
    wire N1075;
    wire N1076;
    wire N1077;
    wire N1078;
    wire N1079;
    wire N1080;
    wire N1081;
    wire N1082;
    wire N1083;
    wire N1084;
    wire N1085;
    wire N1086;
    wire N1087;
    wire N1088;
    wire N1089;
    wire N1090;
    wire N1091;
    wire N1092;
    wire N1093;
    wire N1094;
    wire N1095;
    wire N1096;
    wire N1097;
    wire N1098;
    wire N1099;
    wire N1100;
    wire N1101;
    wire N1102;
    wire N1103;
    wire N1104;
    wire N1105;
    wire N1106;
    wire N1107;
    wire N1108;
    wire N1109;
    wire N1110;
    wire N1111;
    wire N1112;
    wire N1113;
    wire N1114;
    wire N1115;
    wire N1116;
    wire N1117;
    wire N1118;
    wire N1119;
    wire N1120;
    wire N1121;
    wire N1122;
    wire N1123;
    wire N1124;
    wire N1125;
    wire N1126;
    wire N1127;
    wire N1128;
    wire N1129;
    wire N1130;
    wire N1131;
    wire N1132;
    wire N1133;
    wire N1134;
    wire N1135;
    wire N1136;
    wire N1137;
    wire N1138;
    wire N1139;
    wire N1140;
    wire N1141;
    wire N1142;
    wire N1143;
    wire N1144;
    wire N1145;
    wire N1146;
    wire N1147;
    wire N1148;
    wire N1149;
    wire N1150;
    wire N1151;
    wire N1152;
    wire N1153;
    wire N1154;
    wire N1155;
    wire N1156;
    wire N1157;
    wire N1158;
    wire N1159;
    wire N1160;
    wire N1161;
    wire N1162;
    wire N1163;
    wire N1164;
    wire N1165;
    wire N1166;
    wire N1167;
    wire N1168;
    wire N1169;
    wire N1170;
    wire N1171;
    wire N1172;
    wire N1173;
    wire N1174;
    wire N1175;
    wire N1176;
    wire N1177;
    wire N1178;
    wire N1179;
    wire N1180;
    wire N1181;
    wire N1182;
    wire N1183;
    wire N1184;
    wire N1185;
    wire N1186;
    wire N1187;
    wire N1188;
    wire N1189;
    wire N1190;
    wire N1191;
    wire N1192;
    wire N1193;
    wire N1194;
    wire N1195;
    wire N1196;
    wire N1197;
    wire N1198;
    wire N1199;
    wire N1200;
    wire N1201;
    wire N1202;
    wire N1203;
    wire N1204;
    wire N1205;
    wire N1206;
    wire N1207;
    wire N1208;
    wire N1209;
    wire N1210;
    wire N1211;
    wire N1212;
    wire N1213;
    wire N1214;
    wire N1215;
    wire N1216;
    wire N1217;
    wire N1218;
    wire N1219;
    wire N1220;
    wire N1221;
    wire N1222;
    wire N1223;
    wire N1224;
    wire N1225;
    wire N1226;
    wire N1227;
    wire N1228;
    wire N1229;
    wire N1230;
    wire N1231;
    wire N1232;
    wire N1233;
    wire N1234;
    wire N1235;
    wire N1236;
    wire N1237;
    wire N1238;
    wire N1239;
    wire N1240;
    wire N1241;
    wire N1242;
    wire N1243;
    wire N1244;
    wire N1245;
    wire N1246;
    wire N1247;
    wire N1248;
    wire N1249;
    wire N1250;
    wire N1251;
    wire N1252;
    wire N1253;
    wire N1254;
    wire N1255;
    wire N1256;
    wire N1257;
    wire N1258;
    wire N1259;
    wire N1260;
    wire N1261;
    wire N1262;
    wire N1263;
    wire N1264;
    wire N1265;
    wire N1266;
    wire N1267;
    wire N1268;
    wire N1269;
    wire N1270;
    wire N1271;
    wire N1272;
    wire N1273;
    wire N1274;
    wire N1275;
    wire N1276;
    wire N1277;
    wire N1278;
    wire N1279;
    wire N1280;
    wire N1281;
    wire N1282;
    wire N1283;
    wire N1284;
    wire N1285;
    wire N1286;
    wire N1287;
    wire N1288;
    wire N1289;
    wire N1290;
    wire N1291;
    wire N1292;
    wire N1293;
    wire N1294;
    wire N1295;
    wire N1296;
    wire N1297;
    wire N1298;
    wire N1299;
    wire N1300;
    wire N1301;
    wire N1302;
    wire N1303;
    wire N1304;
    wire N1305;
    wire N1306;
    wire N1307;
    wire N1308;
    wire N1309;
    wire N1310;
    wire N1311;
    wire N1312;
    wire N1313;
    wire N1314;
    wire N1315;
    wire N1316;
    wire N1317;
    wire N1318;
    wire N1319;
    wire N1320;
    wire N1321;
    wire N1322;
    wire N1323;
    wire N1324;
    wire N1325;
    wire N1326;
    wire N1327;
    wire N1328;
    wire N1329;
    wire N1330;
    wire N1331;
    wire N1332;
    wire N1333;
    wire N1334;
    wire N1335;
    wire N1336;
    wire N1337;
    wire N1338;
    wire N1339;
    wire N1340;
    wire N1341;
    wire N1342;
    wire N1343;
    wire N1344;
    wire N1345;
    wire N1346;
    wire N1347;
    wire N1348;
    wire N1349;
    wire N1350;
    wire N1351;
    wire N1352;
    wire N1353;
    wire N1354;
    wire N1355;
    wire N1356;
    wire N1357;
    wire N1358;
    wire N1359;
    wire N1360;
    wire N1361;
    wire N1362;
    wire N1363;
    wire N1364;
    wire N1365;
    wire N1366;
    wire N1367;
    wire N1368;
    wire N1369;
    wire N1370;
    wire N1371;
    wire N1372;
    wire N1373;
    wire N1374;
    wire N1375;
    wire N1376;
    wire N1377;
    wire N1378;
    wire N1379;
    wire N1380;
    wire N1381;
    wire N1382;
    wire N1383;
    wire N1384;
    wire N1385;
    wire N1386;
    wire N1387;
    wire N1388;
    wire N1389;
    wire N1390;
    wire N1391;
    wire N1392;
    wire N1393;
    wire N1394;
    wire N1395;
    wire N1396;
    wire N1397;
    wire N1398;
    wire N1399;
    wire N1400;
    wire N1401;
    wire N1402;
    wire N1403;
    wire N1404;
    wire N1405;
    wire N1406;
    wire N1407;
    wire N1408;
    wire N1409;
    wire N1410;
    wire N1411;
    wire N1412;
    wire N1413;
    wire N1414;
    wire N1415;
    wire N1416;
    wire N1417;
    wire N1418;
    wire N1419;
    wire N1420;
    wire N1421;
    wire N1422;
    wire N1423;
    wire N1424;
    wire N1425;
    wire N1426;
    wire N1427;
    wire N1428;
    wire N1429;
    wire N1430;
    wire N1431;
    wire N1432;
    wire N1433;
    wire N1434;
    wire N1435;
    wire N1436;
    wire N1437;
    wire N1438;
    wire N1439;
    wire N1440;
    wire N1441;
    wire N1442;
    wire N1443;
    wire N1444;
    wire N1445;
    wire N1446;
    wire N1447;
    wire N1448;
    wire N1449;
    wire N1450;
    wire N1451;
    wire N1452;
    wire N1453;
    wire N1454;
    wire N1455;
    wire N1456;
    wire N1457;
    wire N1458;
    wire N1459;
    wire N1460;
    wire N1461;
    wire N1462;
    wire N1463;
    wire N1464;
    wire N1465;
    wire N1466;
    wire N1467;
    wire N1468;
    wire N1469;
    wire N1470;
    wire N1471;
    wire N1472;
    wire N1473;
    wire N1474;
    wire N1475;
    wire N1476;
    wire N1477;
    wire N1478;
    wire N1479;
    wire N1480;
    wire N1481;
    wire N1482;
    wire N1483;
    wire N1484;
    wire N1485;
    wire N1486;
    wire N1487;
    wire N1488;
    wire N1489;
    wire N1490;
    wire N1491;
    wire N1492;
    wire N1493;
    wire N1494;
    wire N1495;
    wire N1496;
    wire N1497;
    wire N1498;
    wire N1499;
    wire N1500;
    wire N1501;
    wire N1502;
    wire N1503;
    wire N1504;
    wire N1505;
    wire N1506;
    wire N1507;
    wire N1508;
    wire N1509;
    wire N1510;
    wire N1511;
    wire N1512;
    wire N1513;
    wire N1514;
    wire N1515;
    wire N1516;
    wire N1517;
    wire N1518;
    wire N1519;
    wire N1520;
    wire N1521;
    wire N1522;
    wire N1523;
    wire N1524;
    wire N1525;
    wire N1526;
    wire N1527;
    wire N1528;
    wire N1529;
    wire N1530;
    wire N1531;
    wire N1532;
    wire N1533;
    wire N1534;
    wire N1535;
    wire N1536;
    wire N1537;
    wire N1538;
    wire N1539;
    wire N1540;
    wire N1541;
    wire N1542;
    wire N1543;
    wire N1544;
    wire N1545;
    wire N1546;
    wire N1547;
    wire N1548;
    wire N1549;
    wire N1550;
    wire N1551;
    wire N1552;
    wire N1553;
    wire N1554;
    wire N1555;
    wire N1556;
    wire N1557;
    wire N1558;
    wire N1559;
    wire N1560;
    wire N1561;
    wire N1562;
    wire N1563;
    wire N1564;
    wire N1565;
    wire N1566;
    wire N1567;
    wire N1568;
    wire N1569;
    wire N1570;
    wire N1571;
    wire N1572;
    wire N1573;
    wire N1574;
    wire N1575;
    wire N1576;
    wire N1577;
    wire N1578;
    wire N1579;
    wire N1580;
    wire N1581;
    wire N1582;
    wire N1583;
    wire N1584;
    wire N1585;
    wire N1586;
    wire N1587;
    wire N1588;
    wire N1589;
    wire N1590;
    wire N1591;
    wire N1592;
    wire N1593;
    wire N1594;
    wire N1595;
    wire N1596;
    wire N1597;
    wire N1598;
    wire N1599;
    wire N1600;
    wire N1601;
    wire N1602;
    wire N1603;
    wire N1604;
    wire N1605;
    wire N1606;
    wire N1607;
    wire N1608;
    wire N1609;
    wire N1610;
    wire N1611;
    wire N1612;
    wire N1613;
    wire N1614;
    wire N1615;
    wire N1616;
    wire N1617;
    wire N1618;
    wire N1619;
    wire N1620;
    wire N1621;
    wire N1622;
    wire N1623;
    wire N1624;
    wire N1625;
    wire N1626;
    wire N1627;
    wire N1628;
    wire N1629;
    wire N1630;
    wire N1631;
    wire N1632;
    wire N1633;
    wire N1634;
    wire N1635;
    wire N1636;
    wire N1637;
    wire N1638;
    wire N1639;
    wire N1640;
    wire N1641;
    wire N1642;
    wire N1643;
    wire N1644;
    wire N1645;
    wire N1646;
    wire N1647;
    wire N1648;
    wire N1649;
    wire N1650;
    wire N1651;
    wire N1652;
    wire N1653;
    wire N1654;
    wire N1655;
    wire N1656;
    wire N1657;
    wire N1658;
    wire N1659;
    wire N1660;
    wire N1661;
    wire N1662;
    wire N1663;
    wire N1664;
    wire N1665;
    wire N1666;
    wire N1667;
    wire N1668;
    wire N1669;
    wire N1670;
    wire N1671;
    wire N1672;
    wire N1673;
    wire N1674;
    wire N1675;
    wire N1676;
    wire N1677;
    wire N1678;
    wire N1679;
    wire N1680;
    wire N1681;
    wire N1682;
    wire N1683;
    wire N1684;
    wire N1685;
    wire N1686;
    wire N1687;
    wire N1688;
    wire N1689;
    wire N1690;
    wire N1691;
    wire N1692;
    wire N1693;
    wire N1694;
    wire N1695;
    wire N1696;
    wire N1697;
    wire N1698;
    wire N1699;
    wire N1700;
    wire N1701;
    wire N1702;
    wire N1703;
    wire N1704;
    wire N1705;
    wire N1706;
    wire N1707;
    wire N1708;
    wire N1709;
    wire N1710;
    wire N1711;
    wire N1712;
    wire N1713;
    wire N1714;
    wire N1715;
    wire N1716;
    wire N1717;
    wire N1718;
    wire N1719;
    wire N1720;
    wire N1721;
    wire N1722;
    wire N1723;
    wire N1724;
    wire N1725;
    wire N1726;
    wire N1727;
    wire N1728;
    wire N1729;
    wire N1730;
    wire N1731;
    wire N1732;
    wire N1733;
    wire N1734;
    wire N1735;
    wire N1736;
    wire N1737;
    wire N1738;
    wire N1739;
    wire N1740;
    wire N1741;
    wire N1742;
    wire N1743;
    wire N1744;
    wire N1745;
    wire N1746;
    wire N1747;
    wire N1748;
    wire N1749;
    wire N1750;
    wire N1751;
    wire N1752;
    wire N1753;
    wire N1754;
    wire N1755;
    wire N1756;
    wire N1757;
    wire N1758;
    wire N1759;
    wire N1760;
    wire N1761;
    wire N1762;
    wire N1763;
    wire N1764;
    wire N1765;
    wire N1766;
    wire N1767;
    wire N1768;
    wire N1769;
    wire N1770;
    wire N1771;
    wire N1772;
    wire N1773;
    wire N1774;
    wire N1775;
    wire N1776;
    wire N1777;
    wire N1778;
    wire N1779;
    wire N1780;
    wire N1781;
    wire N1782;
    wire N1783;
    wire N1784;
    wire N1785;
    wire N1786;
    wire N1787;
    wire N1788;
    wire N1789;
    wire N1790;
    wire N1791;
    wire N1792;
    wire N1793;
    wire N1794;
    wire N1795;
    wire N1796;
    wire N1797;
    wire N1798;
    wire N1799;
    wire N1800;
    wire N1801;
    wire N1802;
    wire N1803;
    wire N1804;
    wire N1805;
    wire N1806;
    wire N1807;
    wire N1808;
    wire N1809;
    wire N1810;
    wire N1811;
    wire N1812;
    wire N1813;
    wire N1814;
    wire N1815;
    wire N1816;
    wire N1817;
    wire N1818;
    wire N1819;
    wire N1820;
    wire N1821;
    wire N1822;
    wire N1823;
    wire N1824;
    wire N1825;
    wire N1826;
    wire N1827;
    wire N1828;
    wire N1829;
    wire N1830;
    wire N1831;
    wire N1832;
    wire N1833;
    wire N1834;
    wire N1835;
    wire N1836;
    wire N1837;
    wire N1838;
    wire N1839;
    wire N1840;
    wire N1841;
    wire N1842;
    wire N1843;
    wire N1844;
    wire N1845;
    wire N1846;
    wire N1847;
    wire N1848;
    wire N1849;
    wire N1850;
    wire N1851;
    wire N1852;
    wire N1853;
    wire N1854;
    wire N1855;
    wire N1856;
    wire N1857;
    wire N1858;
    wire N1859;
    wire N1860;
    wire N1861;
    wire N1862;
    wire N1863;
    wire N1864;
    wire N1865;
    wire N1866;
    wire N1867;
    wire N1868;
    wire N1869;
    wire N1870;
    wire N1871;
    wire N1872;
    wire N1873;
    wire N1874;
    wire N1875;
    wire N1876;
    wire N1877;
    wire N1878;
    wire N1879;
    wire N1880;
    wire N1881;
    wire N1882;
    wire N1883;
    wire N1884;
    wire N1885;
    wire N1886;
    wire N1887;
    wire N1888;
    wire N1889;
    wire N1890;
    wire N1891;
    wire N1892;
    wire N1893;
    wire N1894;
    wire N1895;
    wire N1896;
    wire N1897;
    wire N1898;
    wire N1899;
    wire N1900;
    wire N1901;
    wire N1902;
    wire N1903;
    wire N1904;
    wire N1905;
    wire N1906;
    wire N1907;
    wire N1908;
    wire N1909;
    wire N1910;
    wire N1911;
    wire N1912;
    wire N1913;
    wire N1914;
    wire N1915;
    wire N1916;
    wire N1917;
    wire N1918;
    wire N1919;
    wire N1920;
    wire N1921;
    wire N1922;
    wire N1923;
    wire N1924;
    wire N1925;
    wire N1926;
    wire N1927;
    wire N1928;
    wire N1929;
    wire N1930;
    wire N1931;
    wire N1932;
    wire N1933;
    wire N1934;
    wire N1935;
    wire N1936;
    wire N1937;
    wire N1938;
    wire N1939;
    wire N1940;
    wire N1941;
    wire N1942;
    wire N1943;
    wire N1944;
    wire N1945;
    wire N1946;
    wire N1947;
    wire N1948;
    wire N1949;
    wire N1950;
    wire N1951;
    wire N1952;
    wire N1953;
    wire N1954;
    wire N1955;
    wire N1956;
    wire N1957;
    wire N1958;
    wire N1959;
    wire N1960;
    wire N1961;
    wire N1962;
    wire N1963;
    wire N1964;
    wire N1965;
    wire N1966;
    wire N1967;
    wire N1968;
    wire N1969;
    wire N1970;
    wire N1971;
    wire N1972;
    wire N1973;
    wire N1974;
    wire N1975;
    wire N1976;
    wire N1977;
    wire N1978;
    wire N1979;
    wire N1980;
    wire N1981;
    wire N1982;
    wire N1983;
    wire N1984;
    wire N1985;
    wire N1986;
    wire N1987;
    wire N1988;
    wire N1989;
    wire N1990;
    wire N1991;
    wire N1992;
    wire N1993;
    wire N1994;
    wire N1995;
    wire N1996;
    wire N1997;
    wire N1998;
    wire N1999;
    wire N2000;
    wire N2001;
    wire N2002;
    wire N2003;
    wire N2004;
    wire N2005;
    wire N2006;
    wire N2007;
    wire N2008;
    wire N2009;
    wire N2010;
    wire N2011;
    wire N2012;
    wire N2013;
    wire N2014;
    wire N2015;
    wire N2016;
    wire N2017;
    wire N2018;
    wire N2019;
    wire N2020;
    wire N2021;
    wire N2022;
    wire N2023;
    wire N2024;
    wire N2025;
    wire N2026;
    wire N2027;
    wire N2028;
    wire N2029;
    wire N2030;
    wire N2031;
    wire N2032;
    wire N2033;
    wire N2034;
    wire N2035;
    wire N2036;
    wire N2037;
    wire N2038;
    wire N2039;
    wire N2040;
    wire N2041;
    wire N2042;
    wire N2043;
    wire N2044;
    wire N2045;
    wire N2046;
    wire N2047;
    wire N2048;
    wire N2049;
    wire N2050;
    wire N2051;
    wire N2052;
    wire N2053;
    wire N2054;
    wire N2055;
    wire N2056;
    wire N2057;
    wire N2058;
    wire N2059;
    wire N2060;
    wire N2061;
    wire N2062;
    wire N2063;
    wire N2064;
    wire N2065;
    wire N2066;
    wire N2067;
    wire N2068;
    wire N2069;
    wire N2070;
    wire N2071;
    wire N2072;
    wire N2073;
    wire N2074;
    wire N2075;
    wire N2076;
    wire N2077;
    wire N2078;
    wire N2079;
    wire N2080;
    wire N2081;
    wire N2082;
    wire N2083;
    wire N2084;
    wire N2085;
    wire N2086;
    wire N2087;
    wire N2088;
    wire N2089;
    wire N2090;
    wire N2091;
    wire N2092;
    wire N2093;
    wire N2094;
    wire N2095;
    wire N2096;
    wire N2097;
    wire N2098;
    wire N2099;
    wire N2100;
    wire N2101;
    wire N2102;
    wire N2103;
    wire N2104;
    wire N2105;
    wire N2106;
    wire N2107;
    wire N2108;
    wire N2109;
    wire N2110;
    wire N2111;
    wire N2112;
    wire N2113;
    wire N2114;
    wire N2115;
    wire N2116;
    wire N2117;
    wire N2118;
    wire N2119;
    wire N2120;
    wire N2121;
    wire N2122;
    wire N2123;
    wire N2124;
    wire N2125;
    wire N2126;
    wire N2127;
    wire N2128;
    wire N2129;
    wire N2130;
    wire N2131;
    wire N2132;
    wire N2133;
    wire N2134;
    wire N2135;
    wire N2136;
    wire N2137;
    wire N2138;
    wire N2139;
    wire N2140;
    wire N2141;
    wire N2142;
    wire N2143;
    wire N2144;
    wire N2145;
    wire N2146;
    wire N2147;
    wire N2148;
    wire N2149;
    wire N2150;
    wire N2151;
    wire N2152;
    wire N2153;
    wire N2154;
    wire N2155;
    wire N2156;
    wire N2157;
    wire N2158;
    wire N2159;
    wire N2160;
    wire N2161;
    wire N2162;
    wire N2163;
    wire N2164;
    wire N2165;
    wire N2166;
    wire N2167;
    wire N2168;
    wire N2169;
    wire N2170;
    wire N2171;
    wire N2172;
    wire N2173;
    wire N2174;
    wire N2175;
    wire N2176;
    wire N2177;
    wire N2178;
    wire N2179;
    wire N2180;
    wire N2181;
    wire N2182;
    wire N2183;
    wire N2184;
    wire N2185;
    wire N2186;
    wire N2187;
    wire N2188;
    wire N2189;
    wire N2190;
    wire N2191;
    wire N2192;
    wire N2193;
    wire N2194;
    wire N2195;
    wire N2196;
    wire N2197;
    wire N2198;
    wire N2199;
    wire N2200;
    wire N2201;
    wire N2202;
    wire N2203;
    wire N2204;
    wire N2205;
    wire N2206;
    wire N2207;
    wire N2208;
    wire N2209;
    wire N2210;
    wire N2211;
    wire N2212;
    wire N2213;
    wire N2214;
    wire N2215;
    wire N2216;
    wire N2217;
    wire N2218;
    wire N2219;
    wire N2220;
    wire N2221;
    wire N2222;
    wire N2223;
    wire N2224;
    wire N2225;
    wire N2226;
    wire N2227;
    wire N2228;
    wire N2229;
    wire N2230;
    wire N2231;
    wire N2232;
    wire N2233;
    wire N2234;
    wire N2235;
    wire N2236;
    wire N2237;
    wire N2238;
    wire N2239;
    wire N2240;
    wire N2241;
    wire N2242;
    wire N2243;
    wire N2244;
    wire N2245;
    wire N2246;
    wire N2247;
    wire N2248;
    wire N2249;
    wire N2250;
    wire N2251;
    wire N2252;
    wire N2253;
    wire N2254;
    wire N2255;
    wire N2256;
    wire N2257;
    wire N2258;
    wire N2259;
    wire N2260;
    wire N2261;
    wire N2262;
    wire N2263;
    wire N2264;
    wire N2265;
    wire N2266;
    wire N2267;
    wire N2268;
    wire N2269;
    wire N2270;
    wire N2271;
    wire N2272;
    wire N2273;
    wire N2274;
    wire N2275;
    wire N2276;
    wire N2277;
    wire N2278;
    wire N2279;
    wire N2280;
    wire N2281;
    wire N2282;
    wire N2283;
    wire N2284;
    wire N2285;
    wire N2286;
    wire N2287;
    wire N2288;
    wire N2289;
    wire N2290;
    wire N2291;
    wire N2292;
    wire N2293;
    wire N2294;
    wire N2295;
    wire N2296;
    wire N2297;
    wire N2298;
    wire N2299;
    wire N2300;
    wire N2301;
    wire N2302;
    wire N2303;
    wire N2304;
    wire N2305;
    wire N2306;
    wire N2307;
    wire N2308;
    wire N2309;
    wire N2310;
    wire N2311;
    wire N2312;
    wire N2313;
    wire N2314;
    wire N2315;
    wire N2316;
    wire N2317;
    wire N2318;
    wire N2319;
    wire N2320;
    wire N2321;
    wire N2322;
    wire N2323;
    wire N2324;
    wire N2325;
    wire N2326;
    wire N2327;
    wire N2328;
    wire N2329;
    wire N2330;
    wire N2331;
    wire N2332;
    wire N2333;
    wire N2334;
    wire N2335;
    wire N2336;
    wire N2337;
    wire N2338;
    wire N2339;
    wire N2340;
    wire N2341;
    wire N2342;
    wire N2343;
    wire N2344;
    wire N2345;
    wire N2346;
    wire N2347;
    wire N2348;
    wire N2349;
    wire N2350;
    wire N2351;
    wire N2352;
    wire N2353;
    wire N2354;
    wire N2355;
    wire N2356;
    wire N2357;
    wire N2358;
    wire N2359;
    wire N2360;
    wire N2361;
    wire N2362;
    wire N2363;
    wire N2364;
    wire N2365;
    wire N2366;
    wire N2367;
    wire N2368;
    wire N2369;
    wire N2370;
    wire N2371;
    wire N2372;
    wire N2373;
    wire N2374;
    wire N2375;
    wire N2376;
    wire N2377;
    wire N2378;
    wire N2379;
    wire N2380;
    wire N2381;
    wire N2382;
    wire N2383;
    wire N2384;
    wire N2385;
    wire N2386;
    wire N2387;
    wire N2388;
    wire N2389;
    wire N2390;
    wire N2391;
    wire N2392;
    wire N2393;
    wire N2394;
    wire N2395;
    wire N2396;
    wire N2397;
    wire N2398;
    wire N2399;
    wire N2400;
    wire N2401;
    wire N2402;
    wire N2403;
    wire N2404;
    wire N2405;
    wire N2406;
    wire N2407;
    wire N2408;
    wire N2409;
    wire N2410;
    wire N2411;
    wire N2412;
    wire N2413;
    wire N2414;
    wire N2415;
    wire N2416;
    wire N2417;
    wire N2418;
    wire N2419;
    wire N2420;
    wire N2421;
    wire N2422;
    wire N2423;
    wire N2424;
    wire N2425;
    wire N2426;
    wire N2427;
    wire N2428;
    wire N2429;
    wire N2430;
    wire N2431;
    wire N2432;
    wire N2433;
    wire N2434;
    wire N2435;
    wire N2436;
    wire N2437;
    wire N2438;
    wire N2439;
    wire N2440;
    wire N2441;
    wire N2442;
    wire N2443;
    wire N2444;
    wire N2445;
    wire N2446;
    wire N2447;
    wire N2448;
    wire N2449;
    wire N2450;
    wire N2451;
    wire N2452;
    wire N2453;
    wire N2454;
    wire N2455;
    wire N2456;
    wire N2457;
    wire N2458;
    wire N2459;
    wire N2460;
    wire N2461;
    wire N2462;
    wire N2463;
    wire N2464;
    wire N2465;
    wire N2466;
    wire N2467;
    wire N2468;
    wire N2469;
    wire N2470;
    wire N2471;
    wire N2472;
    wire N2473;
    wire N2474;
    wire N2475;
    wire N2476;
    wire N2477;
    wire N2478;
    wire N2479;
    wire N2480;
    wire N2481;
    wire N2482;
    wire N2483;
    wire N2484;
    wire N2485;
    wire N2486;
    wire N2487;
    wire N2488;
    wire N2489;
    wire N2490;
    wire N2491;
    wire N2492;
    wire N2493;
    wire N2494;
    wire N2495;
    wire N2496;
    wire N2497;
    wire N2498;
    wire N2499;
    wire N2500;
    wire N2501;
    wire N2502;
    wire N2503;
    wire N2504;
    wire N2505;
    wire N2506;
    wire N2507;
    wire N2508;
    wire N2509;
    wire N2510;
    wire N2511;
    wire N2512;
    wire N2513;
    wire N2514;
    wire N2515;
    wire N2516;
    wire N2517;
    wire N2518;
    wire N2519;
    wire N2520;
    wire N2521;
    wire N2522;
    wire N2523;
    wire N2524;
    wire N2525;
    wire N2526;
    wire N2527;
    wire N2528;
    wire N2529;
    wire N2530;
    wire N2531;
    wire N2532;
    wire N2533;
    wire N2534;
    wire N2535;
    wire N2536;
    wire N2537;
    wire N2538;
    wire N2539;
    wire N2540;
    wire N2541;
    wire N2542;
    wire N2543;
    wire N2544;
    wire N2545;
    wire N2546;
    wire N2547;
    wire N2548;
    wire N2549;
    wire N2550;
    wire N2551;
    wire N2552;
    wire N2553;
    wire N2554;
    wire N2555;
    wire N2556;
    wire N2557;
    wire N2558;
    wire N2559;
    wire N2560;
    wire N2561;
    wire N2562;
    wire N2563;
    wire N2564;
    wire N2565;
    wire N2566;
    wire N2567;
    wire N2568;
    wire N2569;
    wire N2570;
    wire N2571;
    wire N2572;
    wire N2573;
    wire N2574;
    wire N2575;
    wire N2576;
    wire N2577;
    wire N2578;
    wire N2579;
    wire N2580;
    wire N2581;
    wire N2582;
    wire N2583;
    wire N2584;
    wire N2585;
    wire N2586;
    wire N2587;
    wire N2588;
    wire N2589;
    wire N2590;
    wire N2591;
    wire N2592;
    wire N2593;
    wire N2594;
    wire N2595;
    wire N2596;
    wire N2597;
    wire N2598;
    wire N2599;
    wire N2600;
    wire N2601;
    wire N2602;
    wire N2603;
    wire N2604;
    wire N2605;
    wire N2606;
    wire N2607;
    wire N2608;
    wire N2609;
    wire N2610;
    wire N2611;
    wire N2612;
    wire N2613;
    wire N2614;
    wire N2615;
    wire N2616;
    wire N2617;
    wire N2618;
    wire N2619;
    wire N2620;
    wire N2621;
    wire N2622;
    wire N2623;
    wire N2624;
    wire N2625;
    wire N2626;
    wire N2627;
    wire N2628;
    wire N2629;
    wire N2630;
    wire N2631;
    wire N2632;
    wire N2633;
    wire N2634;
    wire N2635;
    wire N2636;
    wire N2637;
    wire N2638;
    wire N2639;
    wire N2640;
    wire N2641;
    wire N2642;
    wire N2643;
    wire N2644;
    wire N2645;
    wire N2646;
    wire N2647;
    wire N2648;
    wire N2649;
    wire N2650;
    wire N2651;
    wire N2652;
    wire N2653;
    wire N2654;
    wire N2655;
    wire N2656;
    wire N2657;
    wire N2658;
    wire N2659;
    wire N2660;
    wire N2661;
    wire N2662;
    wire N2663;
    wire N2664;
    wire N2665;
    wire N2666;
    wire N2667;
    wire N2668;
    wire N2669;
    wire N2670;
    wire N2671;
    wire N2672;
    wire N2673;
    wire N2674;
    wire N2675;
    wire N2676;
    wire N2677;
    wire N2678;
    wire N2679;
    wire N2680;
    wire N2681;
    wire N2682;
    wire N2683;
    wire N2684;
    wire N2685;
    wire N2686;
    wire N2687;
    wire N2688;
    wire N2689;
    wire N2690;
    wire N2691;
    wire N2692;
    wire N2693;
    wire N2694;
    wire N2695;
    wire N2696;
    wire N2697;
    wire N2698;
    wire N2699;
    wire N2700;
    wire N2701;
    wire N2702;
    wire N2703;
    wire N2704;
    wire N2705;
    wire N2706;
    wire N2707;
    wire N2708;
    wire N2709;
    wire N2710;
    wire N2711;
    wire N2712;
    wire N2713;
    wire N2714;
    wire N2715;
    wire N2716;
    wire N2717;
    wire N2718;
    wire N2719;
    wire N2720;
    wire N2721;
    wire N2722;
    wire N2723;
    wire N2724;
    wire N2725;
    wire N2726;
    wire N2727;
    wire N2728;
    wire N2729;
    wire N2730;
    wire N2731;
    wire N2732;
    wire N2733;
    wire N2734;
    wire N2735;
    wire N2736;
    wire N2737;
    wire N2738;
    wire N2739;
    wire N2740;
    wire N2741;
    wire N2742;
    wire N2743;
    wire N2744;
    wire N2745;
    wire N2746;
    wire N2747;
    wire N2748;
    wire N2749;
    wire N2750;
    wire N2751;
    wire N2752;
    wire N2753;
    wire N2754;
    wire N2755;
    wire N2756;
    wire N2757;
    wire N2758;
    wire N2759;
    wire N2760;
    wire N2761;
    wire N2762;
    wire N2763;
    wire N2764;
    wire N2765;
    wire N2766;
    wire N2767;
    wire N2768;
    wire N2769;
    wire N2770;
    wire N2771;
    wire N2772;
    wire N2773;
    wire N2774;
    wire N2775;
    wire N2776;
    wire N2777;
    wire N2778;
    wire N2779;
    wire N2780;
    wire N2781;
    wire N2782;
    wire N2783;
    wire N2784;
    wire N2785;
    wire N2786;
    wire N2787;
    wire N2788;
    wire N2789;
    wire N2790;
    wire N2791;
    wire N2792;
    wire N2793;
    wire N2794;
    wire N2795;
    wire N2796;
    wire N2797;
    wire N2798;
    wire N2799;
    wire N2800;
    wire N2801;
    wire N2802;
    wire N2803;
    wire N2804;
    wire N2805;
    wire N2806;
    wire N2807;
    wire N2808;
    wire N2809;
    wire N2810;
    wire N2811;
    wire N2812;
    wire N2813;
    wire N2814;
    wire N2815;
    wire N2816;
    wire N2817;
    wire N2818;
    wire N2819;
    wire N2820;
    wire N2821;
    wire N2822;
    wire N2823;
    wire N2824;
    wire N2825;
    wire N2826;
    wire N2827;
    wire N2828;
    wire N2829;
    wire N2830;
    wire N2831;
    wire N2832;
    wire N2833;
    wire N2834;
    wire N2835;
    wire N2836;
    wire N2837;
    wire N2838;
    wire N2839;
    wire N2840;
    wire N2841;
    wire N2842;
    wire N2843;
    wire N2844;
    wire N2845;
    wire N2846;
    wire N2847;
    wire N2848;
    wire N2849;
    wire N2850;
    wire N2851;
    wire N2852;
    wire N2853;
    wire N2854;
    wire N2855;
    wire N2856;
    wire N2857;
    wire N2858;
    wire N2859;
    wire N2860;
    wire N2861;
    wire N2862;
    wire N2863;
    wire N2864;
    wire N2865;
    wire N2866;
    wire N2867;
    wire N2868;
    wire N2869;
    wire N2870;
    wire N2871;
    wire N2872;
    wire N2873;
    wire N2874;
    wire N2875;
    wire N2876;
    wire N2877;
    wire N2878;
    wire N2879;
    wire N2880;
    wire N2881;
    wire N2882;
    wire N2883;
    wire N2884;
    wire N2885;
    wire N2886;
    wire N2887;
    wire N2888;
    wire N2889;
    wire N2890;
    wire N2891;
    wire N2892;
    wire N2893;
    wire N2894;
    wire N2895;
    wire N2896;
    wire N2897;
    wire N2898;
    wire N2899;
    wire N2900;
    wire N2901;
    wire N2902;
    wire N2903;
    wire N2904;
    wire N2905;
    wire N2906;
    wire N2907;
    wire N2908;
    wire N2909;
    wire N2910;
    wire N2911;
    wire N2912;
    wire N2913;
    wire N2914;
    wire N2915;
    wire N2916;
    wire N2917;
    wire N2918;
    wire N2919;
    wire N2920;
    wire N2921;
    wire N2922;
    wire N2923;
    wire N2924;
    wire N2925;
    wire N2926;
    wire N2927;
    wire N2928;
    wire N2929;
    wire N2930;
    wire N2931;
    wire N2932;
    wire N2933;
    wire N2934;
    wire N2935;
    wire N2936;
    wire N2937;
    wire N2938;
    wire N2939;
    wire N2940;
    wire N2941;
    wire N2942;
    wire N2943;
    wire N2944;
    wire N2945;
    wire N2946;
    wire N2947;
    wire N2948;
    wire N2949;
    wire N2950;
    wire N2951;
    wire N2952;
    wire N2953;
    wire N2954;
    wire N2955;
    wire N2956;
    wire N2957;
    wire N2958;
    wire N2959;
    wire N2960;
    wire N2961;
    wire N2962;
    wire N2963;
    wire N2964;
    wire N2965;
    wire N2966;
    wire N2967;
    wire N2968;
    wire N2969;
    wire N2970;
    wire N2971;
    wire N2972;
    wire N2973;
    wire N2974;
    wire N2975;
    wire N2976;
    wire N2977;
    wire N2978;
    wire N2979;
    wire N2980;
    wire N2981;
    wire N2982;
    wire N2983;
    wire N2984;
    wire N2985;
    wire N2986;
    wire N2987;
    wire N2988;
    wire N2989;
    wire N2990;
    wire N2991;
    wire N2992;
    wire N2993;
    wire N2994;
    wire N2995;
    wire N2996;
    wire N2997;
    wire N2998;
    wire N2999;
    wire N3000;
    wire N3001;
    wire N3002;
    wire N3003;
    wire N3004;
    wire N3005;
    wire N3006;
    wire N3007;
    wire N3008;
    wire N3009;
    wire N3010;
    wire N3011;
    wire N3012;
    wire N3013;
    wire N3014;
    wire N3015;
    wire N3016;
    wire N3017;
    wire N3018;
    wire N3019;
    wire N3020;
    wire N3021;
    wire N3022;
    wire N3023;
    wire N3024;
    wire N3025;
    wire N3026;
    wire N3027;
    wire N3028;
    wire N3029;
    wire N3030;
    wire N3031;
    wire N3032;
    wire N3033;
    wire N3034;
    wire N3035;
    wire N3036;
    wire N3037;
    wire N3038;
    wire N3039;
    wire N3040;
    wire N3041;
    wire N3042;
    wire N3043;
    wire N3044;
    wire N3045;
    wire N3046;
    wire N3047;
    wire N3048;
    wire N3049;
    wire N3050;
    wire N3051;
    wire N3052;
    wire N3053;
    wire N3054;
    wire N3055;
    wire N3056;
    wire N3057;
    wire N3058;
    wire N3059;
    wire N3060;
    wire N3061;
    wire N3062;
    wire N3063;
    wire N3064;
    wire N3065;
    wire N3066;
    wire N3067;
    wire N3068;
    wire N3069;
    wire N3070;
    wire N3071;
    wire N3072;
    wire N3073;
    wire N3074;
    wire N3075;
    wire N3076;
    wire N3077;
    wire N3078;
    wire N3079;
    wire N3080;
    wire N3081;
    wire N3082;
    wire N3083;
    wire N3084;
    wire N3085;
    wire N3086;
    wire N3087;
    wire N3088;
    wire N3089;
    wire N3090;
    wire N3091;
    wire N3092;
    wire N3093;
    wire N3094;
    wire N3095;
    wire N3096;
    wire N3097;
    wire N3098;
    wire N3099;
    wire N3100;
    wire N3101;
    wire N3102;
    wire N3103;
    wire N3104;
    wire N3105;
    wire N3106;
    wire N3107;
    wire N3108;
    wire N3109;
    wire N3110;
    wire N3111;
    wire N3112;
    wire N3113;
    wire N3114;
    wire N3115;
    wire N3116;
    wire N3117;
    wire N3118;
    wire N3119;
    wire N3120;
    wire N3121;
    wire N3122;
    wire N3123;
    wire N3124;
    wire N3125;
    wire N3126;
    wire N3127;
    wire N3128;
    wire N3129;
    wire N3130;
    wire N3131;
    wire N3132;
    wire N3133;
    wire N3134;
    wire N3135;
    wire N3136;
    wire N3137;
    wire N3138;
    wire N3139;
    wire N3140;
    wire N3141;
    wire N3142;
    wire N3143;
    wire N3144;
    wire N3145;
    wire N3146;
    wire N3147;
    wire N3148;
    wire N3149;
    wire N3150;
    wire N3151;
    wire N3152;
    wire N3153;
    wire N3154;
    wire N3155;
    wire N3156;
    wire N3157;
    wire N3158;
    wire N3159;
    wire N3160;
    wire N3161;
    wire N3162;
    wire N3163;
    wire N3164;
    wire N3165;
    wire N3166;
    wire N3167;
    wire N3168;
    wire N3169;
    wire N3170;
    wire N3171;
    wire N3172;
    wire N3173;
    wire N3174;
    wire N3175;
    wire N3176;
    wire N3177;
    wire N3178;
    wire N3179;
    wire N3180;
    wire N3181;
    wire N3182;
    wire N3183;
    wire N3184;
    wire N3185;
    wire N3186;
    wire N3187;
    wire N3188;
    wire N3189;
    wire N3190;
    wire N3191;
    wire N3192;
    wire N3193;
    wire N3194;
    wire N3195;
    wire N3196;
    wire N3197;
    wire N3198;
    wire N3199;
    wire N3200;
    wire N3201;
    wire N3202;
    wire N3203;
    wire N3204;
    wire N3205;
    wire N3206;
    wire N3207;
    wire N3208;
    wire N3209;
    wire N3210;
    wire N3211;
    wire N3212;
    wire N3213;
    wire N3214;
    wire N3215;
    wire N3216;
    wire N3217;
    wire N3218;
    wire N3219;
    wire N3220;
    wire N3221;
    wire N3222;
    wire N3223;
    wire N3224;
    wire N3225;
    wire N3226;
    wire N3227;
    wire N3228;
    wire N3229;
    wire N3230;
    wire N3231;
    wire N3232;
    wire N3233;
    wire N3234;
    wire N3235;
    wire N3236;
    wire N3237;
    wire N3238;
    wire N3239;
    wire N3240;
    wire N3241;
    wire N3242;
    wire N3243;
    wire N3244;
    wire N3245;
    wire N3246;
    wire N3247;
    wire N3248;
    wire N3249;
    wire N3250;
    wire N3251;
    wire N3252;
    wire N3253;
    wire N3254;
    wire N3255;
    wire N3256;
    wire N3257;
    wire N3258;
    wire N3259;
    wire N3260;
    wire N3261;
    wire N3262;
    wire N3263;
    wire N3264;
    wire N3265;
    wire N3266;
    wire N3267;
    wire N3268;
    wire N3269;
    wire N3270;
    wire N3271;
    wire N3272;
    wire N3273;
    wire N3274;
    wire N3275;
    wire N3276;
    wire N3277;
    wire N3278;
    wire N3279;
    wire N3280;
    wire N3281;
    wire N3282;
    wire N3283;
    wire N3284;
    wire N3285;
    wire N3286;
    wire N3287;
    wire N3288;
    wire N3289;
    wire N3290;
    wire N3291;
    wire N3292;
    wire N3293;
    wire N3294;
    wire N3295;
    wire N3296;
    wire N3297;
    wire N3298;
    wire N3299;
    wire N3300;
    wire N3301;
    wire N3302;
    wire N3303;
    wire N3304;
    wire N3305;
    wire N3306;
    wire N3307;
    wire N3308;
    wire N3309;
    wire N3310;
    wire N3311;
    wire N3312;
    wire N3313;
    wire N3314;
    wire N3315;
    wire N3316;
    wire N3317;
    wire N3318;
    wire N3319;
    wire N3320;
    wire N3321;
    wire N3322;
    wire N3323;
    wire N3324;
    wire N3325;
    wire N3326;
    wire N3327;
    wire N3328;
    wire N3329;
    wire N3330;
    wire N3331;
    wire N3332;
    wire N3333;
    wire N3334;
    wire N3335;
    wire N3336;
    wire N3337;
    wire N3338;
    wire N3339;
    wire N3340;
    wire N3341;
    wire N3342;
    wire N3343;
    wire N3344;
    wire N3345;
    wire N3346;
    wire N3347;
    wire N3348;
    wire N3349;
    wire N3350;
    wire N3351;
    wire N3352;
    wire N3353;
    wire N3354;
    wire N3355;
    wire N3356;
    wire N3357;
    wire N3358;
    wire N3359;
    wire N3360;
    wire N3361;
    wire N3362;
    wire N3363;
    wire N3364;
    wire N3365;
    wire N3366;
    wire N3367;
    wire N3368;
    wire N3369;
    wire N3370;
    wire N3371;
    wire N3372;
    wire N3373;
    wire N3374;
    wire N3375;
    wire N3376;
    wire N3377;
    wire N3378;
    wire N3379;
    wire N3380;
    wire N3381;
    wire N3382;
    wire N3383;
    wire N3384;
    wire N3385;
    wire N3386;
    wire N3387;
    wire N3388;
    wire N3389;
    wire N3390;
    wire N3391;
    wire N3392;
    wire N3393;
    wire N3394;
    wire N3395;
    wire N3396;
    wire N3397;
    wire N3398;
    wire N3399;
    wire N3400;
    wire N3401;
    wire N3402;
    wire N3403;
    wire N3404;
    wire N3405;
    wire N3406;
    wire N3407;
    wire N3408;
    wire N3409;
    wire N3410;
    wire N3411;
    wire N3412;
    wire N3413;
    wire N3414;
    wire N3415;
    wire N3416;
    wire N3417;
    wire N3418;
    wire N3419;
    wire N3420;
    wire N3421;
    wire N3422;
    wire N3423;
    wire N3424;
    wire N3425;
    wire N3426;
    wire N3427;
    wire N3428;
    wire N3429;
    wire N3430;
    wire N3431;
    wire N3432;
    wire N3433;
    wire N3434;
    wire N3435;
    wire N3436;
    wire N3437;
    wire N3438;
    wire N3439;
    wire N3440;
    wire N3441;
    wire N3442;
    wire N3443;
    wire N3444;
    wire N3445;
    wire N3446;
    wire N3447;
    wire N3448;
    wire N3449;
    wire N3450;
    wire N3451;
    wire N3452;
    wire N3453;
    wire N3454;
    wire N3455;
    wire N3456;
    wire N3457;
    wire N3458;
    wire N3459;
    wire N3460;
    wire N3461;
    wire N3462;
    wire N3463;
    wire N3464;
    wire N3465;
    wire N3466;
    wire N3467;
    wire N3468;
    wire N3469;
    wire N3470;
    wire N3471;
    wire N3472;
    wire N3473;
    wire N3474;
    wire N3475;
    wire N3476;
    wire N3477;
    wire N3478;
    wire N3479;
    wire N3480;
    wire N3481;
    wire N3482;
    wire N3483;
    wire N3484;
    wire N3485;
    wire N3486;
    wire N3487;
    wire N3488;
    wire N3489;
    wire N3490;
    wire N3491;
    wire N3492;
    wire N3493;
    wire N3494;
    wire N3495;
    wire N3496;
    wire N3497;
    wire N3498;
    wire N3499;
    wire N3500;
    wire N3501;
    wire N3502;
    wire N3503;
    wire N3504;
    wire N3505;
    wire N3506;
    wire N3507;
    wire N3508;
    wire N3509;
    wire N3510;
    wire N3511;
    wire N3512;
    wire N3513;
    wire N3514;
    wire N3515;
    wire N3516;
    wire N3517;
    wire N3518;
    wire N3519;
    wire N3520;
    wire N3521;
    wire N3522;
    wire N3523;
    wire N3524;
    wire N3525;
    wire N3526;
    wire N3527;
    wire N3528;
    wire N3529;
    wire N3530;
    wire N3531;
    wire N3532;
    wire N3533;
    wire N3534;
    wire N3535;
    wire N3536;
    wire N3537;
    wire N3538;
    wire N3539;
    wire N3540;
    wire N3541;
    wire N3542;
    wire N3543;
    wire N3544;
    wire N3545;
    wire N3546;
    wire N3547;
    wire N3548;
    wire N3549;
    wire N3550;
    wire N3551;
    wire N3552;
    wire N3553;
    wire N3554;
    wire N3555;
    wire N3556;
    wire N3557;
    wire N3558;
    wire N3559;
    wire N3560;
    wire N3561;
    wire N3562;
    wire N3563;
    wire N3564;
    wire N3565;
    wire N3566;
    wire N3567;
    wire N3568;
    wire N3569;
    wire N3570;
    wire N3571;
    wire N3572;
    wire N3573;
    wire N3574;
    wire N3575;
    wire N3576;
    wire N3577;
    wire N3578;
    wire N3579;
    wire N3580;
    wire N3581;
    wire N3582;
    wire N3583;
    wire N3584;
    wire N3585;
    wire N3586;
    wire N3587;
    wire N3588;
    wire N3589;
    wire N3590;
    wire N3591;
    wire N3592;
    wire N3593;
    wire N3594;
    wire N3595;
    wire N3596;
    wire N3597;
    wire N3598;
    wire N3599;
    wire N3600;
    wire N3601;
    wire N3602;
    wire N3603;
    wire N3604;
    wire N3605;
    wire N3606;
    wire N3607;
    wire N3608;
    wire N3609;
    wire N3610;
    wire N3611;
    wire N3612;
    wire N3613;
    wire N3614;
    wire N3615;
    wire N3616;
    wire N3617;
    wire N3618;
    wire N3619;
    wire N3620;
    wire N3621;
    wire N3622;
    wire N3623;
    wire N3624;
    wire N3625;
    wire N3626;
    wire N3627;
    wire N3628;
    wire N3629;
    wire N3630;
    wire N3631;
    wire N3632;
    wire N3633;
    wire N3634;
    wire N3635;
    wire N3636;
    wire N3637;
    wire N3638;
    wire N3639;
    wire N3640;
    wire N3641;
    wire N3642;
    wire N3643;
    wire N3644;
    wire N3645;
    wire N3646;
    wire N3647;
    wire N3648;
    wire N3649;
    wire N3650;
    wire N3651;
    wire N3652;
    wire N3653;
    wire N3654;
    wire N3655;
    wire N3656;
    wire N3657;
    wire N3658;
    wire N3659;
    wire N3660;
    wire N3661;
    wire N3662;
    wire N3663;
    wire N3664;
    wire N3665;
    wire N3666;
    wire N3667;
    wire N3668;
    wire N3669;
    wire N3670;
    wire N3671;
    wire N3672;
    wire N3673;
    wire N3674;
    wire N3675;
    wire N3676;
    wire N3677;
    wire N3678;
    wire N3679;
    wire N3680;
    wire N3681;
    wire N3682;
    wire N3683;
    wire N3684;
    wire N3685;
    wire N3686;
    wire N3687;
    wire N3688;
    wire N3689;
    wire N3690;
    wire N3691;
    wire N3692;
    wire N3693;
    wire N3694;
    wire N3695;
    wire N3696;
    wire N3697;
    wire N3698;
    wire N3699;
    wire N3700;
    wire N3701;
    wire N3702;
    wire N3703;
    wire N3704;
    wire N3705;
    wire N3706;
    wire N3707;
    wire N3708;
    wire N3709;
    wire N3710;
    wire N3711;
    wire N3712;
    wire N3713;
    wire N3714;
    wire N3715;
    wire N3716;
    wire N3717;
    wire N3718;
    wire N3719;
    wire N3720;
    wire N3721;
    wire N3722;
    wire N3723;
    wire N3724;
    wire N3725;
    wire N3726;
    wire N3727;
    wire N3728;
    wire N3729;
    wire N3730;
    wire N3731;
    wire N3732;
    wire N3733;
    wire N3734;
    wire N3735;
    wire N3736;
    wire N3737;
    wire N3738;
    wire N3739;
    wire N3740;
    wire N3741;
    wire N3742;
    wire N3743;
    wire N3744;
    wire N3745;
    wire N3746;
    wire N3747;
    wire N3748;
    wire N3749;
    wire N3750;
    wire N3751;
    wire N3752;
    wire N3753;
    wire N3754;
    wire N3755;
    wire N3756;
    wire N3757;
    wire N3758;
    wire N3759;
    wire N3760;
    wire N3761;
    wire N3762;
    wire N3763;
    wire N3764;
    wire N3765;
    wire N3766;
    wire N3767;
    wire N3768;
    wire N3769;
    wire N3770;
    wire N3771;
    wire N3772;
    wire N3773;
    wire N3774;
    wire N3775;
    wire N3776;
    wire N3777;
    wire N3778;
    wire N3779;
    wire N3780;
    wire N3781;
    wire N3782;
    wire N3783;
    wire N3784;
    wire N3785;
    wire N3786;
    wire N3787;
    wire N3788;
    wire N3789;
    wire N3790;
    wire N3791;
    wire N3792;
    wire N3793;
    wire N3794;
    wire N3795;
    wire N3796;
    wire N3797;
    wire N3798;
    wire N3799;
    wire N3800;
    wire N3801;
    wire N3802;
    wire N3803;
    wire N3804;
    wire N3805;
    wire N3806;
    wire N3807;
    wire N3808;
    wire N3809;
    wire N3810;
    wire N3811;
    wire N3812;
    wire N3813;
    wire N3814;
    wire N3815;
    wire N3816;
    wire N3817;
    wire N3818;
    wire N3819;
    wire N3820;
    wire N3821;
    wire N3822;
    wire N3823;
    wire N3824;
    wire N3825;
    wire N3826;
    wire N3827;
    wire N3828;
    wire N3829;
    wire N3830;
    wire N3831;
    wire N3832;
    wire N3833;
    wire N3834;
    wire N3835;
    wire N3836;
    wire N3837;
    wire N3838;
    wire N3839;
    wire N3840;
    wire N3841;
    wire N3842;
    wire N3843;
    wire N3844;
    wire N3845;
    wire N3846;
    wire N3847;
    wire N3848;
    wire N3849;
    wire N3850;
    wire N3851;
    wire N3852;
    wire N3853;
    wire N3854;
    wire N3855;
    wire N3856;
    wire N3857;
    wire N3858;
    wire N3859;
    wire N3860;
    wire N3861;
    wire N3862;
    wire N3863;
    wire N3864;
    wire N3865;
    wire N3866;
    wire N3867;
    wire N3868;
    wire N3869;
    wire N3870;
    wire N3871;
    wire N3872;
    wire N3873;
    wire N3874;
    wire N3875;
    wire N3876;
    wire N3877;
    wire N3878;
    wire N3879;
    wire N3880;
    wire N3881;
    wire N3882;
    wire N3883;
    wire N3884;
    wire N3885;
    wire N3886;
    wire N3887;
    wire N3888;
    wire N3889;
    wire N3890;
    wire N3891;
    wire N3892;
    wire N3893;
    wire N3894;
    wire N3895;
    wire N3896;
    wire N3897;
    wire N3898;
    wire N3899;
    wire N3900;
    wire N3901;
    wire N3902;
    wire N3903;
    wire N3904;
    wire N3905;
    wire N3906;
    wire N3907;
    wire N3908;
    wire N3909;
    wire N3910;
    wire N3911;
    wire N3912;
    wire N3913;
    wire N3914;
    wire N3915;
    wire N3916;
    wire N3917;
    wire N3918;
    wire N3919;
    wire N3920;
    wire N3921;
    wire N3922;
    wire N3923;
    wire N3924;
    wire N3925;
    wire N3926;
    wire N3927;
    wire N3928;
    wire N3929;
    wire N3930;
    wire N3931;
    wire N3932;
    wire N3933;
    wire N3934;
    wire N3935;
    wire N3936;
    wire N3937;
    wire N3938;
    wire N3939;
    wire N3940;
    wire N3941;
    wire N3942;
    wire N3943;
    wire N3944;
    wire N3945;
    wire N3946;
	INVX1 g_N386 (N215, N386);
	INVX1 g_N387 (N1045, N387);
	AND2X1 g_N388 (N2519, N2678, N388);
	BUFX2 g_N389 (N3530, N389);
	INVX1 g_N390 (N1592, N390);
	BUFX2 g_N391 (N1399, N391);
	BUFX2 g_N392 (N3538, N392);
	INVX1 g_N393 (N1691, N393);
	INVX1 g_N394 (N1169, N394);
	INVX1 g_N395 (N3353, N395);
	BUFX2 g_N396 (N3623, N396);
	INVX1 g_N397 (N2570, N397);
	AND2X1 g_N398 (N1998, N1149, N398);
	AND2X1 g_N399 (N1213, N2886, N399);
	BUFX2 g_N400 (N3287, N400);
	AND2X1 g_N401 (N3009, N2791, N401);
	AND2X1 g_N402 (N1731, N1171, N402);
	INVX1 g_N403 (N2926, N403);
	BUFX2 g_N404 (N1783, N404);
	AND2X1 g_N405 (N1786, N1554, N405);
	AND2X1 g_N406 (N3358, N416, N406);
	INVX1 g_N407 (N3838, N407);
	BUFX2 g_N257 (N1379, N257);
	BUFX2 g_N408 (N2731, N408);
	BUFX2 g_N409 (N3224, N409);
	BUFX2 g_N410 (N2263, N410);
	INVX1 g_N411 (N2784, N411);
	AND2X1 g_N412 (N3756, N3587, N412);
	INVX1 g_N413 (N3447, N413);
	INVX1 g_N414 (N2960, N414);
	INVX1 g_N415 (N981, N415);
	INVX1 g_N416 (N2131, N416);
	AND2X1 g_N417 (N621, N3441, N417);
	INVX1 g_N418 (N3078, N418);
	INVX1 g_N419 (N65, N419);
	INVX1 g_N420 (N855, N420);
	INVX1 g_N421 (N185, N421);
	INVX1 g_N422 (N841, N422);
	INVX1 g_N423 (N558, N423);
	AND2X1 g_N424 (N1508, N1797, N424);
	BUFX2 g_N425 (N1222, N425);
	INVX1 g_N426 (N187, N426);
	AND2X1 g_N427 (N3047, N3048, N427);
	INVX1 g_N428 (N1992, N428);
	INVX1 g_N429 (N147, N429);
	INVX1 g_N430 (N168, N430);
	INVX1 g_N431 (N1154, N431);
	INVX1 g_N432 (N1470, N432);
	BUFX2 g_N433 (N3187, N433);
	INVX1 g_N434 (N1513, N434);
	AND2X1 g_N435 (N3784, N2250, N435);
	INVX1 g_N436 (N1293, N436);
	BUFX2 g_N437 (N2370, N437);
	INVX1 g_N438 (N2285, N438);
	BUFX2 g_N439 (N2417, N439);
	AND2X1 g_N440 (N3600, N2381, N440);
	AND2X1 g_N441 (N1534, N2253, N441);
	INVX1 g_N442 (N3793, N442);
	BUFX2 g_N443 (N509, N443);
	BUFX2 g_N444 (N3180, N444);
	BUFX2 g_N445 (N1026, N445);
	INVX1 g_N446 (N1500, N446);
	INVX1 g_N447 (N2858, N447);
	INVX1 g_N448 (N1790, N448);
	AND2X1 g_N449 (N256, N147, N449);
	BUFX2 g_N450 (N3826, N450);
	INVX1 g_N451 (N251, N451);
	INVX1 g_N452 (N496, N452);
	INVX1 g_N453 (N1683, N453);
	BUFX2 g_N454 (N1516, N454);
	BUFX2 g_N455 (N2437, N455);
	AND2X1 g_N456 (N3554, N3610, N456);
	BUFX2 g_N457 (N1268, N457);
	BUFX2 g_N458 (N3565, N458);
	BUFX2 g_N459 (N2907, N459);
	INVX1 g_N460 (N210, N460);
	INVX1 g_N461 (N554, N461);
	BUFX2 g_N462 (N449, N462);
	BUFX2 g_N463 (N1936, N463);
	BUFX2 g_N464 (N586, N464);
	INVX1 g_N465 (N2381, N465);
	BUFX2 g_N466 (N2147, N466);
	AND2X1 g_N467 (N895, N1089, N467);
	INVX1 g_N468 (N2331, N468);
	AND2X1 g_N469 (N3093, N2668, N469);
	INVX1 g_N470 (N162, N470);
	INVX1 g_N471 (N2834, N471);
	INVX1 g_N472 (N583, N472);
	BUFX2 g_N473 (N2796, N473);
	BUFX2 g_N474 (N1288, N474);
	BUFX2 g_N475 (N3785, N475);
	BUFX2 g_N476 (N3718, N476);
	AND2X1 g_N477 (N1427, N1116, N477);
	INVX1 g_N478 (N55, N478);
	BUFX2 g_N479 (N2982, N479);
	BUFX2 g_N258 (N3304, N258);
	AND2X1 g_N480 (N1255, N3439, N480);
	BUFX2 g_N481 (N1538, N481);
	INVX1 g_N482 (N9, N482);
	BUFX2 g_N483 (N2161, N483);
	INVX1 g_N484 (N566, N484);
	AND2X1 g_N485 (N2048, N2910, N485);
	AND2X1 g_N486 (N3400, N414, N486);
	BUFX2 g_N487 (N848, N487);
	INVX1 g_N488 (N223, N488);
	AND2X1 g_N489 (N432, N1083, N489);
	AND2X1 g_N490 (N1198, N687, N490);
	INVX1 g_N491 (N2848, N491);
	INVX1 g_N492 (N3751, N492);
	AND2X1 g_N493 (N471, N2158, N493);
	BUFX2 g_N494 (N3936, N494);
	INVX1 g_N495 (N2149, N495);
	BUFX2 g_N496 (N1165, N496);
	AND2X1 g_N497 (N2927, N1995, N497);
	INVX1 g_N498 (N130, N498);
	BUFX2 g_N499 (N3199, N499);
	BUFX2 g_N500 (N3408, N500);
	BUFX2 g_N501 (N935, N501);
	INVX1 g_N502 (N3837, N502);
	BUFX2 g_N503 (N2934, N503);
	INVX1 g_N504 (N175, N504);
	BUFX2 g_N259 (N1759, N259);
	AND2X1 g_N505 (N420, N3503, N505);
	INVX1 g_N506 (N3746, N506);
	INVX1 g_N507 (N2137, N507);
	BUFX2 g_N508 (N497, N508);
	AND2X1 g_N509 (N3742, N1956, N509);
	AND2X1 g_N510 (N2086, N2104, N510);
	INVX1 g_N511 (N3531, N511);
	INVX1 g_N512 (N3854, N512);
	INVX1 g_N513 (N92, N513);
	AND2X1 g_N514 (N1042, N1911, N514);
	INVX1 g_N515 (N2699, N515);
	INVX1 g_N516 (N540, N516);
	INVX1 g_N517 (N1849, N517);
	BUFX2 g_N518 (N1640, N518);
	AND2X1 g_N519 (N2473, N2969, N519);
	BUFX2 g_N520 (N1705, N520);
	INVX1 g_N521 (N455, N521);
	BUFX2 g_N522 (N3096, N522);
	BUFX2 g_N523 (N1775, N523);
	BUFX2 g_N524 (N705, N524);
	INVX1 g_N525 (N212, N525);
	INVX1 g_N526 (N3196, N526);
	AND2X1 g_N527 (N48, N1, N527);
	AND2X1 g_N528 (N2464, N1254, N528);
	INVX1 g_N529 (N2088, N529);
	AND2X1 g_N530 (N1745, N2711, N530);
	INVX1 g_N531 (N1195, N531);
	INVX1 g_N532 (N145, N532);
	INVX1 g_N533 (N2636, N533);
	BUFX2 g_N534 (N1425, N534);
	INVX1 g_N535 (N1161, N535);
	INVX1 g_N536 (N189, N536);
	BUFX2 g_N537 (N857, N537);
	INVX1 g_N538 (N2661, N538);
	BUFX2 g_N539 (N3707, N539);
	BUFX2 g_N540 (N528, N540);
	BUFX2 g_N541 (N1559, N541);
	INVX1 g_N542 (N2689, N542);
	AND2X1 g_N543 (N1921, N2973, N543);
	AND2X1 g_N544 (N2958, N964, N544);
	BUFX2 g_N545 (N1857, N545);
	BUFX2 g_N546 (N435, N546);
	INVX1 g_N547 (N3385, N547);
	INVX1 g_N548 (N2743, N548);
	INVX1 g_N549 (N1485, N549);
	BUFX2 g_N550 (N2344, N550);
	INVX1 g_N551 (N2494, N551);
	INVX1 g_N552 (N2329, N552);
	BUFX2 g_N260 (N466, N260);
	INVX1 g_N553 (N3277, N553);
	BUFX2 g_N554 (N562, N554);
	BUFX2 g_N261 (N3033, N261);
	INVX1 g_N555 (N105, N555);
	AND2X1 g_N556 (N2562, N2007, N556);
	AND2X1 g_N557 (N619, N1829, N557);
	BUFX2 g_N558 (N3567, N558);
	BUFX2 g_N559 (N3845, N559);
	INVX1 g_N560 (N2520, N560);
	AND2X1 g_N561 (N2512, N470, N561);
	AND2X1 g_N562 (N3617, N478, N562);
	INVX1 g_N563 (N1660, N563);
	INVX1 g_N564 (N1957, N564);
	INVX1 g_N565 (N404, N565);
	BUFX2 g_N566 (N3121, N566);
	INVX1 g_N567 (N2576, N567);
	AND2X1 g_N568 (N960, N957, N568);
	INVX1 g_N569 (N3864, N569);
	BUFX2 g_N570 (N868, N570);
	INVX1 g_N571 (N3886, N571);
	BUFX2 g_N572 (N3637, N572);
	BUFX2 g_N262 (N2408, N262);
	BUFX2 g_N573 (N1152, N573);
	BUFX2 g_N574 (N1002, N574);
	INVX1 g_N575 (N102, N575);
	INVX1 g_N576 (N2295, N576);
	AND2X1 g_N577 (N3384, N2980, N577);
	BUFX2 g_N578 (N2998, N578);
	AND2X1 g_N579 (N2042, N533, N579);
	BUFX2 g_N580 (N3873, N580);
	INVX1 g_N581 (N1502, N581);
	BUFX2 g_N582 (N3661, N582);
	BUFX2 g_N583 (N947, N583);
	INVX1 g_N584 (N3037, N584);
	INVX1 g_N585 (N2067, N585);
	AND2X1 g_N586 (N395, N2833, N586);
	AND2X1 g_N587 (N887, N3550, N587);
	AND2X1 g_N588 (N134, N161, N588);
	BUFX2 g_N589 (N3155, N589);
	INVX1 g_N590 (N3940, N590);
	INVX1 g_N591 (N1895, N591);
	AND2X1 g_N592 (N3015, N2761, N592);
	INVX1 g_N593 (N3902, N593);
	AND2X1 g_N594 (N2243, N448, N594);
	BUFX2 g_N595 (N2455, N595);
	BUFX2 g_N596 (N1150, N596);
	INVX1 g_N597 (N255, N597);
	INVX1 g_N598 (N153, N598);
	BUFX2 g_N263 (N2767, N263);
	BUFX2 g_N599 (N3703, N599);
	AND2X1 g_N600 (N2544, N2577, N600);
	BUFX2 g_N264 (N473, N264);
	BUFX2 g_N601 (N771, N601);
	INVX1 g_N602 (N3054, N602);
	AND2X1 g_N603 (N2171, N2505, N603);
	AND2X1 g_N604 (N691, N891, N604);
	INVX1 g_N605 (N128, N605);
	AND2X1 g_N606 (N3183, N2616, N606);
	BUFX2 g_N265 (N3580, N265);
	INVX1 g_N607 (N2976, N607);
	AND2X1 g_N608 (N133, N187, N608);
	AND2X1 g_N609 (N28, N102, N609);
	AND2X1 g_N610 (N984, N3644, N610);
	INVX1 g_N611 (N3628, N611);
	AND2X1 g_N612 (N430, N3666, N612);
	AND2X1 g_N613 (N3040, N2402, N613);
	INVX1 g_N614 (N151, N614);
	BUFX2 g_N615 (N1280, N615);
	BUFX2 g_N266 (N2380, N266);
	INVX1 g_N616 (N3335, N616);
	BUFX2 g_N617 (N3773, N617);
	BUFX2 g_N618 (N1654, N618);
	INVX1 g_N619 (N2384, N619);
	INVX1 g_N620 (N731, N620);
	INVX1 g_N621 (N50, N621);
	BUFX2 g_N622 (N3822, N622);
	INVX1 g_N623 (N97, N623);
	AND2X1 g_N624 (N791, N1104, N624);
	BUFX2 g_N625 (N1865, N625);
	AND2X1 g_N626 (N3612, N2075, N626);
	INVX1 g_N627 (N1400, N627);
	BUFX2 g_N628 (N1853, N628);
	INVX1 g_N629 (N26, N629);
	AND2X1 g_N630 (N896, N2955, N630);
	INVX1 g_N631 (N1167, N631);
	AND2X1 g_N632 (N1217, N1791, N632);
	INVX1 g_N633 (N445, N633);
	INVX1 g_N634 (N1195, N634);
	AND2X1 g_N635 (N2291, N1943, N635);
	BUFX2 g_N636 (N2382, N636);
	BUFX2 g_N637 (N3698, N637);
	BUFX2 g_N638 (N1476, N638);
	BUFX2 g_N639 (N1690, N639);
	AND2X1 g_N640 (N1825, N1754, N640);
	AND2X1 g_N641 (N3783, N3394, N641);
	BUFX2 g_N642 (N3930, N642);
	AND2X1 g_N643 (N3432, N2483, N643);
	INVX1 g_N644 (N524, N644);
	BUFX2 g_N645 (N2052, N645);
	BUFX2 g_N646 (N3852, N646);
	INVX1 g_N647 (N1491, N647);
	INVX1 g_N648 (N905, N648);
	BUFX2 g_N649 (N2239, N649);
	AND2X1 g_N650 (N2385, N2552, N650);
	AND2X1 g_N651 (N1411, N3748, N651);
	INVX1 g_N652 (N596, N652);
	BUFX2 g_N653 (N1539, N653);
	BUFX2 g_N654 (N3167, N654);
	AND2X1 g_N655 (N923, N507, N655);
	INVX1 g_N656 (N2492, N656);
	BUFX2 g_N657 (N2467, N657);
	AND2X1 g_N658 (N1472, N521, N658);
	BUFX2 g_N659 (N816, N659);
	AND2X1 g_N660 (N2679, N3171, N660);
	AND2X1 g_N661 (N894, N933, N661);
	BUFX2 g_N662 (N878, N662);
	BUFX2 g_N663 (N2947, N663);
	INVX1 g_N664 (N163, N664);
	INVX1 g_N665 (N1024, N665);
	BUFX2 g_N666 (N3527, N666);
	BUFX2 g_N667 (N2363, N667);
	INVX1 g_N668 (N1622, N668);
	INVX1 g_N669 (N813, N669);
	BUFX2 g_N670 (N3865, N670);
	AND2X1 g_N671 (N2594, N1897, N671);
	INVX1 g_N672 (N599, N672);
	AND2X1 g_N673 (N2999, N2895, N673);
	BUFX2 g_N674 (N1912, N674);
	BUFX2 g_N675 (N3473, N675);
	AND2X1 g_N676 (N3045, N2922, N676);
	BUFX2 g_N677 (N2566, N677);
	BUFX2 g_N678 (N1518, N678);
	INVX1 g_N679 (N3348, N679);
	AND2X1 g_N680 (N2040, N2556, N680);
	AND2X1 g_N681 (N859, N457, N681);
	BUFX2 g_N682 (N3943, N682);
	BUFX2 g_N267 (N885, N267);
	BUFX2 g_N268 (N2813, N268);
	INVX1 g_N683 (N1358, N683);
	INVX1 g_N684 (N2156, N684);
	INVX1 g_N685 (N1258, N685);
	AND2X1 g_N686 (N86, N222, N686);
	INVX1 g_N687 (N2065, N687);
	INVX1 g_N688 (N2493, N688);
	BUFX2 g_N689 (N2632, N689);
	BUFX2 g_N690 (N2421, N690);
	INVX1 g_N691 (N3037, N691);
	INVX1 g_N692 (N101, N692);
	INVX1 g_N693 (N3492, N693);
	AND2X1 g_N694 (N2332, N1210, N694);
	AND2X1 g_N695 (N1503, N988, N695);
	INVX1 g_N696 (N1526, N696);
	INVX1 g_N697 (N3782, N697);
	AND2X1 g_N698 (N97, N51, N698);
	BUFX2 g_N699 (N2841, N699);
	INVX1 g_N700 (N2172, N700);
	INVX1 g_N701 (N574, N701);
	INVX1 g_N702 (N3361, N702);
	BUFX2 g_N703 (N1846, N703);
	AND2X1 g_N704 (N1703, N1190, N704);
	AND2X1 g_N705 (N442, N3855, N705);
	INVX1 g_N706 (N880, N706);
	AND2X1 g_N707 (N3125, N452, N707);
	INVX1 g_N708 (N1478, N708);
	AND2X1 g_N709 (N789, N3570, N709);
	AND2X1 g_N710 (N1738, N2793, N710);
	BUFX2 g_N711 (N658, N711);
	AND2X1 g_N712 (N3298, N3896, N712);
	BUFX2 g_N713 (N2502, N713);
	AND2X1 g_N714 (N167, N206, N714);
	AND2X1 g_N715 (N3348, N3363, N715);
	INVX1 g_N716 (N2848, N716);
	BUFX2 g_N717 (N783, N717);
	INVX1 g_N718 (N2441, N718);
	INVX1 g_N719 (N3710, N719);
	INVX1 g_N720 (N204, N720);
	INVX1 g_N721 (N86, N721);
	INVX1 g_N722 (N3899, N722);
	INVX1 g_N723 (N3254, N723);
	BUFX2 g_N724 (N920, N724);
	INVX1 g_N725 (N3280, N725);
	INVX1 g_N726 (N3129, N726);
	BUFX2 g_N269 (N1905, N269);
	AND2X1 g_N727 (N3510, N1406, N727);
	AND2X1 g_N728 (N2744, N2056, N728);
	AND2X1 g_N729 (N428, N564, N729);
	BUFX2 g_N730 (N2655, N730);
	BUFX2 g_N731 (N1270, N731);
	AND2X1 g_N732 (N2520, N526, N732);
	AND2X1 g_N733 (N2904, N623, N733);
	AND2X1 g_N734 (N3000, N788, N734);
	INVX1 g_N735 (N850, N735);
	AND2X1 g_N736 (N1450, N1659, N736);
	AND2X1 g_N737 (N3729, N3124, N737);
	BUFX2 g_N738 (N1537, N738);
	BUFX2 g_N739 (N2915, N739);
	INVX1 g_N740 (N2378, N740);
	INVX1 g_N741 (N2393, N741);
	AND2X1 g_N742 (N3014, N2708, N742);
	INVX1 g_N743 (N2433, N743);
	AND2X1 g_N744 (N18, N163, N744);
	INVX1 g_N745 (N3489, N745);
	BUFX2 g_N746 (N2728, N746);
	BUFX2 g_N747 (N3605, N747);
	INVX1 g_N748 (N667, N748);
	INVX1 g_N749 (N841, N749);
	INVX1 g_N750 (N68, N750);
	BUFX2 g_N751 (N1646, N751);
	INVX1 g_N752 (N67, N752);
	INVX1 g_N753 (N445, N753);
	BUFX2 g_N270 (N1704, N270);
	AND2X1 g_N754 (N2735, N1084, N754);
	INVX1 g_N755 (N206, N755);
	AND2X1 g_N756 (N970, N1075, N756);
	INVX1 g_N757 (N2506, N757);
	BUFX2 g_N758 (N3120, N758);
	AND2X1 g_N759 (N2619, N2759, N759);
	BUFX2 g_N760 (N3480, N760);
	AND2X1 g_N761 (N2510, N1756, N761);
	INVX1 g_N762 (N3350, N762);
	INVX1 g_N763 (N3559, N763);
	BUFX2 g_N764 (N2885, N764);
	INVX1 g_N765 (N2216, N765);
	INVX1 g_N766 (N1902, N766);
	INVX1 g_N767 (N856, N767);
	INVX1 g_N768 (N1372, N768);
	INVX1 g_N769 (N636, N769);
	AND2X1 g_N770 (N855, N3469, N770);
	AND2X1 g_N771 (N538, N3062, N771);
	BUFX2 g_N271 (N2701, N271);
	AND2X1 g_N772 (N1064, N1828, N772);
	BUFX2 g_N773 (N2693, N773);
	AND2X1 g_N774 (N3680, N1076, N774);
	AND2X1 g_N775 (N2893, N749, N775);
	BUFX2 g_N776 (N1051, N776);
	AND2X1 g_N777 (N1632, N1656, N777);
	BUFX2 g_N778 (N977, N778);
	INVX1 g_N779 (N2609, N779);
	AND2X1 g_N780 (N2586, N3022, N780);
	BUFX2 g_N781 (N1658, N781);
	INVX1 g_N782 (N618, N782);
	AND2X1 g_N783 (N2801, N633, N783);
	INVX1 g_N784 (N2318, N784);
	AND2X1 g_N785 (N2090, N958, N785);
	AND2X1 g_N786 (N917, N2091, N786);
	AND2X1 g_N787 (N1931, N1058, N787);
	INVX1 g_N788 (N747, N788);
	INVX1 g_N789 (N108, N789);
	INVX1 g_N790 (N1144, N790);
	INVX1 g_N791 (N3764, N791);
	INVX1 g_N792 (N1540, N792);
	INVX1 g_N793 (N14, N793);
	AND2X1 g_N794 (N2315, N1109, N794);
	INVX1 g_N795 (N2144, N795);
	BUFX2 g_N796 (N1688, N796);
	INVX1 g_N797 (N213, N797);
	BUFX2 g_N798 (N1722, N798);
	INVX1 g_N799 (N2404, N799);
	AND2X1 g_N800 (N2994, N3501, N800);
	INVX1 g_N801 (N1374, N801);
	AND2X1 g_N802 (N1079, N2584, N802);
	AND2X1 g_N803 (N3311, N2613, N803);
	INVX1 g_N804 (N2850, N804);
	BUFX2 g_N805 (N1296, N805);
	INVX1 g_N806 (N1240, N806);
	AND2X1 g_N807 (N1834, N1603, N807);
	INVX1 g_N808 (N96, N808);
	AND2X1 g_N809 (N2851, N996, N809);
	BUFX2 g_N810 (N3027, N810);
	AND2X1 g_N811 (N585, N975, N811);
	INVX1 g_N812 (N3059, N812);
	BUFX2 g_N813 (N955, N813);
	INVX1 g_N814 (N3110, N814);
	BUFX2 g_N815 (N2669, N815);
	AND2X1 g_N816 (N3024, N1586, N816);
	AND2X1 g_N817 (N189, N232, N817);
	BUFX2 g_N818 (N3847, N818);
	AND2X1 g_N819 (N2968, N1536, N819);
	BUFX2 g_N820 (N2423, N820);
	BUFX2 g_N821 (N1715, N821);
	AND2X1 g_N822 (N2034, N801, N822);
	INVX1 g_N823 (N1549, N823);
	BUFX2 g_N824 (N2762, N824);
	INVX1 g_N825 (N1189, N825);
	AND2X1 g_N826 (N1021, N397, N826);
	BUFX2 g_N827 (N2564, N827);
	INVX1 g_N828 (N1263, N828);
	INVX1 g_N829 (N1129, N829);
	INVX1 g_N830 (N3594, N830);
	INVX1 g_N831 (N3150, N831);
	INVX1 g_N832 (N3432, N832);
	AND2X1 g_N833 (N3160, N647, N833);
	AND2X1 g_N834 (N426, N1289, N834);
	BUFX2 g_N835 (N707, N835);
	INVX1 g_N836 (N37, N836);
	INVX1 g_N837 (N3903, N837);
	BUFX2 g_N838 (N3247, N838);
	INVX1 g_N839 (N43, N839);
	INVX1 g_N840 (N3672, N840);
	BUFX2 g_N841 (N2269, N841);
	AND2X1 g_N842 (N910, N1147, N842);
	INVX1 g_N843 (N2045, N843);
	AND2X1 g_N844 (N34, N74, N844);
	AND2X1 g_N845 (N3005, N3486, N845);
	BUFX2 g_N272 (N3505, N272);
	BUFX2 g_N273 (N3728, N273);
	BUFX2 g_N846 (N655, N846);
	BUFX2 g_N847 (N1716, N847);
	AND2X1 g_N848 (N2089, N1692, N848);
	INVX1 g_N849 (N670, N849);
	BUFX2 g_N850 (N3722, N850);
	AND2X1 g_N851 (N1025, N2311, N851);
	INVX1 g_N852 (N3793, N852);
	AND2X1 g_N853 (N752, N3179, N853);
	AND2X1 g_N854 (N506, N1158, N854);
	BUFX2 g_N855 (N3534, N855);
	BUFX2 g_N856 (N3257, N856);
	AND2X1 g_N857 (N3290, N2357, N857);
	AND2X1 g_N858 (N512, N1066, N858);
	INVX1 g_N859 (N3211, N859);
	AND2X1 g_N860 (N921, N3905, N860);
	AND2X1 g_N861 (N852, N2222, N861);
	BUFX2 g_N862 (N3914, N862);
	AND2X1 g_N863 (N77, N162, N863);
	INVX1 g_N864 (N1819, N864);
	INVX1 g_N865 (N98, N865);
	AND2X1 g_N866 (N3803, N3932, N866);
	AND2X1 g_N867 (N142, N11, N867);
	AND2X1 g_N868 (N2462, N1769, N868);
	AND2X1 g_N869 (N1711, N3426, N869);
	BUFX2 g_N870 (N3662, N870);
	INVX1 g_N871 (N2501, N871);
	INVX1 g_N872 (N83, N872);
	INVX1 g_N873 (N197, N873);
	INVX1 g_N874 (N2644, N874);
	BUFX2 g_N274 (N3882, N274);
	BUFX2 g_N875 (N3115, N875);
	INVX1 g_N876 (N2754, N876);
	INVX1 g_N877 (N207, N877);
	AND2X1 g_N878 (N1350, N652, N878);
	BUFX2 g_N879 (N2188, N879);
	BUFX2 g_N880 (N3416, N880);
	INVX1 g_N881 (N678, N881);
	AND2X1 g_N882 (N622, N415, N882);
	AND2X1 g_N883 (N2084, N1464, N883);
	BUFX2 g_N884 (N985, N884);
	BUFX2 g_N885 (N2901, N885);
	INVX1 g_N886 (N1022, N886);
	INVX1 g_N887 (N2314, N887);
	BUFX2 g_N888 (N2125, N888);
	BUFX2 g_N889 (N834, N889);
	BUFX2 g_N890 (N1836, N890);
	BUFX2 g_N891 (N2412, N891);
	AND2X1 g_N892 (N2574, N1947, N892);
	BUFX2 g_N893 (N1256, N893);
	INVX1 g_N894 (N410, N894);
	INVX1 g_N895 (N3864, N895);
	INVX1 g_N896 (N731, N896);
	AND2X1 g_N897 (N3226, N1847, N897);
	AND2X1 g_N898 (N1781, N1415, N898);
	INVX1 g_N899 (N2806, N899);
	BUFX2 g_N900 (N2717, N900);
	INVX1 g_N901 (N1975, N901);
	BUFX2 g_N902 (N2705, N902);
	AND2X1 g_N903 (N3518, N1040, N903);
	BUFX2 g_N904 (N1497, N904);
	BUFX2 g_N905 (N2231, N905);
	AND2X1 g_N906 (N3581, N2630, N906);
	BUFX2 g_N907 (N2478, N907);
	AND2X1 g_N908 (N1707, N3808, N908);
	INVX1 g_N909 (N3918, N909);
	BUFX2 g_N910 (N1523, N910);
	BUFX2 g_N911 (N2607, N911);
	BUFX2 g_N912 (N3790, N912);
	INVX1 g_N913 (N1863, N913);
	BUFX2 g_N914 (N715, N914);
	INVX1 g_N915 (N3834, N915);
	INVX1 g_N916 (N3082, N916);
	INVX1 g_N917 (N200, N917);
	INVX1 g_N918 (N250, N918);
	BUFX2 g_N275 (N1391, N275);
	BUFX2 g_N919 (N1133, N919);
	AND2X1 g_N920 (N2406, N1854, N920);
	BUFX2 g_N921 (N1474, N921);
	BUFX2 g_N922 (N2168, N922);
	INVX1 g_N923 (N921, N923);
	INVX1 g_N924 (N3946, N924);
	AND2X1 g_N925 (N75, N79, N925);
	INVX1 g_N926 (N1415, N926);
	BUFX2 g_N927 (N3860, N927);
	INVX1 g_N928 (N2391, N928);
	BUFX2 g_N929 (N1942, N929);
	BUFX2 g_N930 (N1266, N930);
	BUFX2 g_N931 (N3456, N931);
	AND2X1 g_N932 (N2888, N1070, N932);
	INVX1 g_N933 (N3721, N933);
	INVX1 g_N934 (N2310, N934);
	AND2X1 g_N935 (N104, N250, N935);
	INVX1 g_N936 (N900, N936);
	AND2X1 g_N937 (N991, N1893, N937);
	AND2X1 g_N938 (N3815, N2152, N938);
	AND2X1 g_N939 (N3274, N3248, N939);
	AND2X1 g_N940 (N209, N98, N940);
	BUFX2 g_N941 (N3392, N941);
	INVX1 g_N942 (N3712, N942);
	INVX1 g_N943 (N3129, N943);
	INVX1 g_N944 (N2249, N944);
	BUFX2 g_N945 (N3245, N945);
	AND2X1 g_N946 (N2839, N3275, N946);
	AND2X1 g_N947 (N3866, N2978, N947);
	AND2X1 g_N948 (N3201, N963, N948);
	INVX1 g_N949 (N2650, N949);
	INVX1 g_N950 (N1616, N950);
	AND2X1 g_N951 (N2025, N2983, N951);
	AND2X1 g_N952 (N3111, N3598, N952);
	BUFX2 g_N953 (N1841, N953);
	BUFX2 g_N954 (N2602, N954);
	AND2X1 g_N955 (N2124, N3491, N955);
	INVX1 g_N956 (N1030, N956);
	INVX1 g_N957 (N2170, N957);
	BUFX2 g_N958 (N946, N958);
	AND2X1 g_N959 (N81, N179, N959);
	INVX1 g_N960 (N396, N960);
	BUFX2 g_N961 (N2822, N961);
	AND2X1 g_N962 (N516, N2954, N962);
	BUFX2 g_N963 (N2919, N963);
	INVX1 g_N964 (N2032, N964);
	BUFX2 g_N276 (N2647, N276);
	BUFX2 g_N965 (N2143, N965);
	BUFX2 g_N966 (N2734, N966);
	BUFX2 g_N967 (N2292, N967);
	BUFX2 g_N277 (N2811, N277);
	INVX1 g_N968 (N2992, N968);
	INVX1 g_N969 (N1899, N969);
	INVX1 g_N970 (N1219, N970);
	INVX1 g_N971 (N3502, N971);
	BUFX2 g_N972 (N1229, N972);
	AND2X1 g_N973 (N2255, N982, N973);
	AND2X1 g_N974 (N3762, N840, N974);
	INVX1 g_N975 (N617, N975);
	BUFX2 g_N976 (N2815, N976);
	AND2X1 g_N977 (N3736, N3031, N977);
	INVX1 g_N978 (N3346, N978);
	AND2X1 g_N979 (N3092, N1844, N979);
	INVX1 g_N980 (N2007, N980);
	BUFX2 g_N981 (N3455, N981);
	INVX1 g_N982 (N181, N982);
	INVX1 g_N983 (N1957, N983);
	INVX1 g_N984 (N2232, N984);
	AND2X1 g_N985 (N2166, N3305, N985);
	AND2X1 g_N986 (N1301, N3630, N986);
	BUFX2 g_N987 (N1446, N987);
	INVX1 g_N988 (N573, N988);
	INVX1 g_N989 (N2049, N989);
	AND2X1 g_N990 (N3163, N2404, N990);
	INVX1 g_N991 (N165, N991);
	INVX1 g_N992 (N2781, N992);
	INVX1 g_N993 (N1246, N993);
	INVX1 g_N994 (N475, N994);
	INVX1 g_N995 (N3011, N995);
	INVX1 g_N996 (N1327, N996);
	BUFX2 g_N997 (N613, N997);
	INVX1 g_N998 (N2939, N998);
	AND2X1 g_N999 (N2288, N3454, N999);
	AND2X1 g_N1000 (N1232, N2022, N1000);
	INVX1 g_N1001 (N545, N1001);
	AND2X1 g_N1002 (N2083, N1793, N1002);
	BUFX2 g_N1003 (N3026, N1003);
	AND2X1 g_N1004 (N2772, N743, N1004);
	AND2X1 g_N1005 (N130, N136, N1005);
	BUFX2 g_N278 (N3003, N278);
	BUFX2 g_N1006 (N579, N1006);
	BUFX2 g_N1007 (N2130, N1007);
	INVX1 g_N1008 (N2331, N1008);
	INVX1 g_N1009 (N1597, N1009);
	BUFX2 g_N1010 (N3759, N1010);
	INVX1 g_N1011 (N2501, N1011);
	AND2X1 g_N1012 (N13, N178, N1012);
	BUFX2 g_N1013 (N2557, N1013);
	BUFX2 g_N1014 (N467, N1014);
	INVX1 g_N1015 (N1790, N1015);
	INVX1 g_N1016 (N682, N1016);
	INVX1 g_N1017 (N474, N1017);
	INVX1 g_N1018 (N10, N1018);
	AND2X1 g_N1019 (N2534, N2517, N1019);
	INVX1 g_N1020 (N927, N1020);
	INVX1 g_N1021 (N3492, N1021);
	BUFX2 g_N1022 (N1582, N1022);
	BUFX2 g_N1023 (N3182, N1023);
	BUFX2 g_N1024 (N1481, N1024);
	INVX1 g_N1025 (N45, N1025);
	AND2X1 g_N1026 (N1315, N750, N1026);
	BUFX2 g_N1027 (N1153, N1027);
	AND2X1 g_N1028 (N174, N202, N1028);
	AND2X1 g_N1029 (N3877, N1733, N1029);
	BUFX2 g_N1030 (N2077, N1030);
	INVX1 g_N1031 (N929, N1031);
	AND2X1 g_N1032 (N3596, N3839, N1032);
	BUFX2 g_N1033 (N505, N1033);
	INVX1 g_N1034 (N2642, N1034);
	INVX1 g_N1035 (N3, N1035);
	AND2X1 g_N1036 (N1579, N1227, N1036);
	AND2X1 g_N1037 (N2857, N3519, N1037);
	AND2X1 g_N1038 (N1514, N2260, N1038);
	BUFX2 g_N1039 (N2027, N1039);
	INVX1 g_N1040 (N225, N1040);
	BUFX2 g_N1041 (N2853, N1041);
	INVX1 g_N1042 (N3902, N1042);
	INVX1 g_N1043 (N238, N1043);
	BUFX2 g_N1044 (N3085, N1044);
	BUFX2 g_N1045 (N424, N1045);
	BUFX2 g_N1046 (N3517, N1046);
	BUFX2 g_N1047 (N3122, N1047);
	BUFX2 g_N1048 (N1816, N1048);
	INVX1 g_N1049 (N1880, N1049);
	INVX1 g_N1050 (N22, N1050);
	AND2X1 g_N1051 (N1747, N1668, N1051);
	INVX1 g_N1052 (N2259, N1052);
	AND2X1 g_N1053 (N943, N2030, N1053);
	AND2X1 g_N1054 (N2558, N3074, N1054);
	BUFX2 g_N1055 (N1319, N1055);
	AND2X1 g_N1056 (N790, N1606, N1056);
	BUFX2 g_N1057 (N1220, N1057);
	INVX1 g_N1058 (N1944, N1058);
	INVX1 g_N1059 (N3858, N1059);
	INVX1 g_N1060 (N3211, N1060);
	AND2X1 g_N1061 (N1566, N2210, N1061);
	BUFX2 g_N1062 (N427, N1062);
	BUFX2 g_N1063 (N3468, N1063);
	INVX1 g_N1064 (N2914, N1064);
	AND2X1 g_N1065 (N1691, N1442, N1065);
	INVX1 g_N1066 (N1980, N1066);
	BUFX2 g_N1067 (N882, N1067);
	AND2X1 g_N1068 (N2783, N1533, N1068);
	INVX1 g_N1069 (N625, N1069);
	BUFX2 g_N1070 (N2185, N1070);
	BUFX2 g_N1071 (N809, N1071);
	AND2X1 g_N1072 (N971, N2294, N1072);
	AND2X1 g_N1073 (N2424, N2524, N1073);
	BUFX2 g_N1074 (N587, N1074);
	INVX1 g_N1075 (N1486, N1075);
	INVX1 g_N1076 (N911, N1076);
	BUFX2 g_N1077 (N3843, N1077);
	INVX1 g_N1078 (N3634, N1078);
	INVX1 g_N1079 (N123, N1079);
	AND2X1 g_N1080 (N2348, N2784, N1080);
	BUFX2 g_N1081 (N3170, N1081);
	BUFX2 g_N1082 (N802, N1082);
	BUFX2 g_N1083 (N3547, N1083);
	BUFX2 g_N1084 (N2070, N1084);
	BUFX2 g_N1085 (N2173, N1085);
	BUFX2 g_N1086 (N681, N1086);
	INVX1 g_N1087 (N1529, N1087);
	INVX1 g_N1088 (N2473, N1088);
	INVX1 g_N1089 (N677, N1089);
	BUFX2 g_N1090 (N2537, N1090);
	INVX1 g_N1091 (N2224, N1091);
	INVX1 g_N1092 (N2503, N1092);
	INVX1 g_N1093 (N2251, N1093);
	INVX1 g_N1094 (N2241, N1094);
	AND2X1 g_N1095 (N1720, N503, N1095);
	INVX1 g_N1096 (N1466, N1096);
	AND2X1 g_N1097 (N2737, N2804, N1097);
	INVX1 g_N1098 (N3884, N1098);
	INVX1 g_N1099 (N3503, N1099);
	INVX1 g_N1100 (N2749, N1100);
	INVX1 g_N1101 (N1611, N1101);
	INVX1 g_N1102 (N2927, N1102);
	BUFX2 g_N279 (N3738, N279);
	BUFX2 g_N280 (N730, N280);
	INVX1 g_N1103 (N539, N1103);
	INVX1 g_N1104 (N1923, N1104);
	INVX1 g_N1105 (N1572, N1105);
	AND2X1 g_N1106 (N1059, N1676, N1106);
	BUFX2 g_N1107 (N770, N1107);
	INVX1 g_N1108 (N3713, N1108);
	INVX1 g_N1109 (N3348, N1109);
	AND2X1 g_N1110 (N1748, N1101, N1110);
	INVX1 g_N1111 (N617, N1111);
	BUFX2 g_N1112 (N2600, N1112);
	INVX1 g_N1113 (N3080, N1113);
	INVX1 g_N1114 (N194, N1114);
	AND2X1 g_N1115 (N1859, N768, N1115);
	INVX1 g_N1116 (N3389, N1116);
	AND2X1 g_N1117 (N198, N230, N1117);
	AND2X1 g_N1118 (N3628, N2189, N1118);
	BUFX2 g_N1119 (N2755, N1119);
	INVX1 g_N1120 (N208, N1120);
	AND2X1 g_N1121 (N1488, N1099, N1121);
	AND2X1 g_N1122 (N3664, N3326, N1122);
	AND2X1 g_N1123 (N190, N14, N1123);
	AND2X1 g_N1124 (N3478, N3771, N1124);
	AND2X1 g_N1125 (N1827, N2428, N1125);
	INVX1 g_N1126 (N1210, N1126);
	BUFX2 g_N1127 (N908, N1127);
	INVX1 g_N1128 (N572, N1128);
	BUFX2 g_N1129 (N1584, N1129);
	INVX1 g_N1130 (N1413, N1130);
	INVX1 g_N1131 (N2756, N1131);
	AND2X1 g_N1132 (N2559, N1611, N1132);
	AND2X1 g_N1133 (N3229, N2812, N1133);
	BUFX2 g_N1134 (N1525, N1134);
	AND2X1 g_N1135 (N3747, N1458, N1135);
	AND2X1 g_N1136 (N3039, N2942, N1136);
	INVX1 g_N1137 (N2374, N1137);
	AND2X1 g_N1138 (N1193, N2471, N1138);
	AND2X1 g_N1139 (N235, N58, N1139);
	BUFX2 g_N1140 (N1810, N1140);
	INVX1 g_N1141 (N3069, N1141);
	INVX1 g_N1142 (N2924, N1142);
	AND2X1 g_N1143 (N740, N2542, N1143);
	BUFX2 g_N1144 (N3727, N1144);
	AND2X1 g_N1145 (N238, N78, N1145);
	BUFX2 g_N1146 (N2780, N1146);
	INVX1 g_N1147 (N1505, N1147);
	INVX1 g_N1148 (N2413, N1148);
	INVX1 g_N1149 (N3409, N1149);
	AND2X1 g_N1150 (N1287, N3195, N1150);
	AND2X1 g_N1151 (N1882, N909, N1151);
	AND2X1 g_N1152 (N3211, N1892, N1152);
	AND2X1 g_N1153 (N3232, N3236, N1153);
	BUFX2 g_N1154 (N1344, N1154);
	INVX1 g_N1155 (N1261, N1155);
	AND2X1 g_N1156 (N2064, N3406, N1156);
	INVX1 g_N1157 (N1400, N1157);
	INVX1 g_N1158 (N3254, N1158);
	AND2X1 g_N1159 (N3430, N1812, N1159);
	INVX1 g_N1160 (N254, N1160);
	BUFX2 g_N281 (N3057, N281);
	BUFX2 g_N1161 (N600, N1161);
	AND2X1 g_N1162 (N2527, N2816, N1162);
	INVX1 g_N1163 (N1140, N1163);
	BUFX2 g_N282 (N1175, N282);
	INVX1 g_N1164 (N3915, N1164);
	AND2X1 g_N1165 (N149, N215, N1165);
	AND2X1 g_N1166 (N994, N3917, N1166);
	BUFX2 g_N1167 (N2732, N1167);
	BUFX2 g_N1168 (N1320, N1168);
	BUFX2 g_N1169 (N2683, N1169);
	BUFX2 g_N1170 (N1917, N1170);
	INVX1 g_N1171 (N2952, N1171);
	AND2X1 g_N1172 (N2252, N1700, N1172);
	INVX1 g_N1173 (N3110, N1173);
	BUFX2 g_N1174 (N510, N1174);
	BUFX2 g_N1175 (N869, N1175);
	BUFX2 g_N1176 (N2496, N1176);
	INVX1 g_N1177 (N2258, N1177);
	BUFX2 g_N1178 (N2150, N1178);
	INVX1 g_N1179 (N891, N1179);
	INVX1 g_N1180 (N3649, N1180);
	BUFX2 g_N1181 (N3923, N1181);
	AND2X1 g_N1182 (N1424, N2293, N1182);
	INVX1 g_N1183 (N2051, N1183);
	AND2X1 g_N1184 (N2541, N2044, N1184);
	INVX1 g_N1185 (N1920, N1185);
	AND2X1 g_N1186 (N122, N192, N1186);
	AND2X1 g_N1187 (N3300, N836, N1187);
	INVX1 g_N1188 (N2922, N1188);
	BUFX2 g_N1189 (N3227, N1189);
	INVX1 g_N1190 (N1335, N1190);
	INVX1 g_N1191 (N80, N1191);
	AND2X1 g_N1192 (N194, N140, N1192);
	INVX1 g_N1193 (N3892, N1193);
	BUFX2 g_N1194 (N1843, N1194);
	BUFX2 g_N1195 (N3352, N1195);
	INVX1 g_N1196 (N249, N1196);
	AND2X1 g_N1197 (N3431, N1573, N1197);
	INVX1 g_N1198 (N3190, N1198);
	INVX1 g_N1199 (N1146, N1199);
	BUFX2 g_N1200 (N3006, N1200);
	AND2X1 g_N1201 (N3381, N2720, N1201);
	INVX1 g_N1202 (N1880, N1202);
	INVX1 g_N1203 (N1430, N1203);
	BUFX2 g_N283 (N2675, N283);
	INVX1 g_N1204 (N1602, N1204);
	AND2X1 g_N1205 (N1396, N2060, N1205);
	INVX1 g_N1206 (N900, N1206);
	INVX1 g_N1207 (N1849, N1207);
	AND2X1 g_N1208 (N247, N211, N1208);
	BUFX2 g_N284 (N1346, N284);
	AND2X1 g_N1209 (N1403, N835, N1209);
	BUFX2 g_N1210 (N2575, N1210);
	INVX1 g_N1211 (N1862, N1211);
	INVX1 g_N1212 (N601, N1212);
	INVX1 g_N1213 (N2050, N1213);
	AND2X1 g_N1214 (N1910, N2704, N1214);
	AND2X1 g_N1215 (N847, N1866, N1215);
	INVX1 g_N1216 (N2429, N1216);
	INVX1 g_N1217 (N3647, N1217);
	BUFX2 g_N1218 (N1870, N1218);
	BUFX2 g_N1219 (N3331, N1219);
	AND2X1 g_N1220 (N2439, N918, N1220);
	BUFX2 g_N1221 (N1591, N1221);
	AND2X1 g_N1222 (N3346, N3590, N1222);
	INVX1 g_N1223 (N1259, N1223);
	BUFX2 g_N1224 (N1028, N1224);
	AND2X1 g_N1225 (N1204, N1617, N1225);
	INVX1 g_N1226 (N3143, N1226);
	INVX1 g_N1227 (N2300, N1227);
	BUFX2 g_N1228 (N1005, N1228);
	AND2X1 g_N1229 (N3102, N3438, N1229);
	INVX1 g_N1230 (N3093, N1230);
	AND2X1 g_N1231 (N3868, N3579, N1231);
	INVX1 g_N1232 (N115, N1232);
	INVX1 g_N1233 (N1014, N1233);
	AND2X1 g_N1234 (N76, N216, N1234);
	BUFX2 g_N1235 (N3881, N1235);
	AND2X1 g_N1236 (N1609, N3603, N1236);
	BUFX2 g_N1237 (N1357, N1237);
	INVX1 g_N1238 (N66, N1238);
	AND2X1 g_N1239 (N484, N3811, N1239);
	BUFX2 g_N1240 (N1056, N1240);
	BUFX2 g_N1241 (N3083, N1241);
	INVX1 g_N1242 (N2489, N1242);
	AND2X1 g_N1243 (N1365, N2035, N1243);
	INVX1 g_N1244 (N1926, N1244);
	AND2X1 g_N1245 (N3629, N3786, N1245);
	BUFX2 g_N1246 (N1187, N1246);
	AND2X1 g_N1247 (N1307, N1423, N1247);
	INVX1 g_N1248 (N167, N1248);
	AND2X1 g_N1249 (N1351, N907, N1249);
	INVX1 g_N1250 (N1806, N1250);
	INVX1 g_N1251 (N3564, N1251);
	BUFX2 g_N1252 (N543, N1252);
	AND2X1 g_N1253 (N249, N3682, N1253);
	INVX1 g_N1254 (N1877, N1254);
	INVX1 g_N1255 (N2195, N1255);
	AND2X1 g_N1256 (N3752, N876, N1256);
	BUFX2 g_N1257 (N490, N1257);
	BUFX2 g_N1258 (N1727, N1258);
	BUFX2 g_N1259 (N2963, N1259);
	BUFX2 g_N1260 (N469, N1260);
	BUFX2 g_N1261 (N3551, N1261);
	INVX1 g_N1262 (N1510, N1262);
	BUFX2 g_N1263 (N952, N1263);
	AND2X1 g_N1264 (N1230, N1168, N1264);
	BUFX2 g_N1265 (N486, N1265);
	AND2X1 g_N1266 (N877, N1160, N1266);
	INVX1 g_N1267 (N1398, N1267);
	AND2X1 g_N1268 (N2965, N3329, N1268);
	INVX1 g_N1269 (N835, N1269);
	AND2X1 g_N1270 (N125, N217, N1270);
	INVX1 g_N1271 (N1590, N1271);
	BUFX2 g_N1272 (N3133, N1272);
	AND2X1 g_N1273 (N1269, N436, N1273);
	INVX1 g_N1274 (N3386, N1274);
	INVX1 g_N1275 (N890, N1275);
	AND2X1 g_N1276 (N109, N67, N1276);
	AND2X1 g_N1277 (N1034, N2099, N1277);
	BUFX2 g_N1278 (N1205, N1278);
	INVX1 g_N1279 (N3337, N1279);
	AND2X1 g_N1280 (N3599, N3219, N1280);
	INVX1 g_N1281 (N2162, N1281);
	INVX1 g_N1282 (N2368, N1282);
	INVX1 g_N1283 (N3272, N1283);
	INVX1 g_N1284 (N1944, N1284);
	INVX1 g_N1285 (N921, N1285);
	INVX1 g_N1286 (N3800, N1286);
	INVX1 g_N1287 (N3302, N1287);
	AND2X1 g_N1288 (N899, N461, N1288);
	INVX1 g_N1289 (N133, N1289);
	INVX1 g_N1290 (N1920, N1290);
	BUFX2 g_N1291 (N2010, N1291);
	AND2X1 g_N1292 (N2664, N1521, N1292);
	BUFX2 g_N1293 (N1839, N1293);
	INVX1 g_N1294 (N2889, N1294);
	BUFX2 g_N1295 (N787, N1295);
	AND2X1 g_N1296 (N784, N2775, N1296);
	AND2X1 g_N1297 (N1670, N3325, N1297);
	INVX1 g_N1298 (N3627, N1298);
	AND2X1 g_N1299 (N1216, N511, N1299);
	AND2X1 g_N1300 (N2470, N2395, N1300);
	INVX1 g_N1301 (N1127, N1301);
	BUFX2 g_N1302 (N2721, N1302);
	INVX1 g_N1303 (N3540, N1303);
	BUFX2 g_N285 (N3376, N285);
	INVX1 g_N1304 (N252, N1304);
	AND2X1 g_N1305 (N2550, N3658, N1305);
	BUFX2 g_N286 (N3802, N286);
	INVX1 g_N1306 (N2427, N1306);
	INVX1 g_N1307 (N1698, N1307);
	AND2X1 g_N1308 (N224, N151, N1308);
	AND2X1 g_N1309 (N3659, N3850, N1309);
	BUFX2 g_N1310 (N1277, N1310);
	AND2X1 g_N1311 (N1303, N1970, N1311);
	BUFX2 g_N1312 (N1249, N1312);
	BUFX2 g_N1313 (N2148, N1313);
	BUFX2 g_N1314 (N1845, N1314);
	INVX1 g_N1315 (N160, N1315);
	AND2X1 g_N1316 (N779, N1281, N1316);
	BUFX2 g_N1317 (N3690, N1317);
	BUFX2 g_N1318 (N632, N1318);
	AND2X1 g_N1319 (N2304, N2076, N1319);
	AND2X1 g_N1320 (N3388, N1020, N1320);
	AND2X1 g_N1321 (N2625, N3589, N1321);
	BUFX2 g_N287 (N3070, N287);
	BUFX2 g_N1322 (N2880, N1322);
	AND2X1 g_N1323 (N525, N2618, N1323);
	AND2X1 g_N1324 (N3944, N3020, N1324);
	AND2X1 g_N1325 (N3848, N3267, N1325);
	BUFX2 g_N1326 (N530, N1326);
	BUFX2 g_N1327 (N2624, N1327);
	BUFX2 g_N1328 (N2548, N1328);
	BUFX2 g_N1329 (N3307, N1329);
	INVX1 g_N1330 (N2309, N1330);
	INVX1 g_N1331 (N954, N1331);
	AND2X1 g_N1332 (N248, N73, N1332);
	BUFX2 g_N1333 (N2452, N1333);
	INVX1 g_N1334 (N1486, N1334);
	BUFX2 g_N1335 (N2826, N1335);
	INVX1 g_N1336 (N558, N1336);
	INVX1 g_N1337 (N2806, N1337);
	BUFX2 g_N1338 (N1695, N1338);
	AND2X1 g_N1339 (N3136, N2274, N1339);
	BUFX2 g_N1340 (N3911, N1340);
	INVX1 g_N1341 (N2248, N1341);
	BUFX2 g_N288 (N537, N288);
	BUFX2 g_N1342 (N732, N1342);
	BUFX2 g_N1343 (N786, N1343);
	AND2X1 g_N1344 (N3146, N1183, N1344);
	INVX1 g_N1345 (N987, N1345);
	BUFX2 g_N1346 (N568, N1346);
	INVX1 g_N1347 (N2660, N1347);
	AND2X1 g_N1348 (N146, N20, N1348);
	INVX1 g_N1349 (N1318, N1349);
	INVX1 g_N1350 (N2845, N1350);
	INVX1 g_N1351 (N2200, N1351);
	AND2X1 g_N1352 (N3440, N3626, N1352);
	AND2X1 g_N1353 (N152, N24, N1353);
	BUFX2 g_N1354 (N2114, N1354);
	AND2X1 g_N1355 (N92, N84, N1355);
	INVX1 g_N1356 (N1477, N1356);
	AND2X1 g_N1357 (N3434, N551, N1357);
	BUFX2 g_N1358 (N733, N1358);
	AND2X1 g_N1359 (N234, N129, N1359);
	AND2X1 g_N1360 (N1991, N3772, N1360);
	AND2X1 g_N1361 (N741, N2312, N1361);
	INVX1 g_N1362 (N2565, N1362);
	INVX1 g_N1363 (N99, N1363);
	INVX1 g_N1364 (N1318, N1364);
	INVX1 g_N1365 (N3350, N1365);
	AND2X1 g_N1366 (N1948, N1027, N1366);
	INVX1 g_N1367 (N487, N1367);
	AND2X1 g_N1368 (N2017, N1400, N1368);
	AND2X1 g_N1369 (N812, N3872, N1369);
	INVX1 g_N1370 (N1809, N1370);
	AND2X1 g_N1371 (N634, N1557, N1371);
	BUFX2 g_N1372 (N1073, N1372);
	AND2X1 g_N1373 (N3906, N563, N1373);
	BUFX2 g_N1374 (N3487, N1374);
	BUFX2 g_N1375 (N1225, N1375);
	INVX1 g_N1376 (N1246, N1376);
	INVX1 g_N1377 (N2509, N1377);
	INVX1 g_N1378 (N1709, N1378);
	BUFX2 g_N1379 (N3382, N1379);
	BUFX2 g_N289 (N3428, N289);
	AND2X1 g_N1380 (N1437, N3184, N1380);
	AND2X1 g_N1381 (N3508, N2159, N1381);
	INVX1 g_N1382 (N3478, N1382);
	AND2X1 g_N1383 (N3148, N584, N1383);
	INVX1 g_N1384 (N2939, N1384);
	BUFX2 g_N1385 (N3754, N1385);
	AND2X1 g_N1386 (N3410, N3814, N1386);
	AND2X1 g_N1387 (N2179, N1011, N1387);
	INVX1 g_N1388 (N3524, N1388);
	INVX1 g_N1389 (N3595, N1389);
	INVX1 g_N1390 (N2032, N1390);
	BUFX2 g_N1391 (N2760, N1391);
	INVX1 g_N1392 (N1826, N1392);
	AND2X1 g_N1393 (N1069, N1016, N1393);
	INVX1 g_N1394 (N3511, N1394);
	BUFX2 g_N1395 (N1780, N1395);
	INVX1 g_N1396 (N3368, N1396);
	INVX1 g_N1397 (N81, N1397);
	BUFX2 g_N1398 (N1624, N1398);
	AND2X1 g_N1399 (N2773, N721, N1399);
	BUFX2 g_N1400 (N1758, N1400);
	AND2X1 g_N1401 (N875, N2648, N1401);
	BUFX2 g_N1402 (N1479, N1402);
	INVX1 g_N1403 (N2510, N1403);
	BUFX2 g_N1404 (N1097, N1404);
	INVX1 g_N1405 (N2599, N1405);
	INVX1 g_N1406 (N2200, N1406);
	BUFX2 g_N1407 (N2750, N1407);
	INVX1 g_N1408 (N3466, N1408);
	BUFX2 g_N1409 (N3017, N1409);
	BUFX2 g_N1410 (N671, N1410);
	INVX1 g_N1411 (N158, N1411);
	AND2X1 g_N1412 (N1284, N2913, N1412);
	BUFX2 g_N1413 (N1901, N1413);
	AND2X1 g_N1414 (N1142, N3775, N1414);
	BUFX2 g_N1415 (N1757, N1415);
	BUFX2 g_N1416 (N2190, N1416);
	BUFX2 g_N1417 (N2896, N1417);
	INVX1 g_N1418 (N3613, N1418);
	AND2X1 g_N1419 (N2299, N1494, N1419);
	INVX1 g_N1420 (N907, N1420);
	INVX1 g_N1421 (N38, N1421);
	INVX1 g_N1422 (N2926, N1422);
	INVX1 g_N1423 (N1683, N1423);
	INVX1 g_N1424 (N3668, N1424);
	AND2X1 g_N1425 (N128, N126, N1425);
	AND2X1 g_N1426 (N3153, N1444, N1426);
	BUFX2 g_N1427 (N3123, N1427);
	BUFX2 g_N1428 (N2449, N1428);
	BUFX2 g_N1429 (N2268, N1429);
	BUFX2 g_N1430 (N937, N1430);
	BUFX2 g_N1431 (N1728, N1431);
	INVX1 g_N1432 (N541, N1432);
	INVX1 g_N1433 (N3715, N1433);
	AND2X1 g_N1434 (N239, N54, N1434);
	BUFX2 g_N1435 (N1509, N1435);
	AND2X1 g_N1436 (N3507, N482, N1436);
	INVX1 g_N1437 (N143, N1437);
	AND2X1 g_N1438 (N3555, N3296, N1438);
	AND2X1 g_N1439 (N3940, N2254, N1439);
	BUFX2 g_N1440 (N1612, N1440);
	BUFX2 g_N1441 (N2867, N1441);
	BUFX2 g_N290 (N3700, N290);
	INVX1 g_N1442 (N3470, N1442);
	AND2X1 g_N1443 (N1851, N1111, N1443);
	INVX1 g_N1444 (N2295, N1444);
	INVX1 g_N1445 (N3819, N1445);
	AND2X1 g_N1446 (N2436, N2908, N1446);
	AND2X1 g_N1447 (N1623, N3281, N1447);
	BUFX2 g_N1448 (N2906, N1448);
	BUFX2 g_N1449 (N1490, N1449);
	BUFX2 g_N1450 (N2047, N1450);
	INVX1 g_N1451 (N244, N1451);
	BUFX2 g_N1452 (N1192, N1452);
	AND2X1 g_N1453 (N61, N171, N1453);
	INVX1 g_N1454 (N1260, N1454);
	AND2X1 g_N1455 (N2686, N3713, N1455);
	INVX1 g_N1456 (N1964, N1456);
	INVX1 g_N1457 (N1697, N1457);
	INVX1 g_N1458 (N820, N1458);
	INVX1 g_N1459 (N3223, N1459);
	INVX1 g_N1460 (N890, N1460);
	AND2X1 g_N1461 (N1663, N1639, N1461);
	AND2X1 g_N1462 (N1768, N2515, N1462);
	AND2X1 g_N1463 (N3648, N2764, N1463);
	INVX1 g_N1464 (N1129, N1464);
	BUFX2 g_N1465 (N694, N1465);
	BUFX2 g_N1466 (N527, N1466);
	BUFX2 g_N1467 (N2580, N1467);
	BUFX2 g_N1468 (N1940, N1468);
	AND2X1 g_N1469 (N389, N2990, N1469);
	BUFX2 g_N1470 (N3706, N1470);
	INVX1 g_N1471 (N2834, N1471);
	INVX1 g_N1472 (N1717, N1472);
	INVX1 g_N1473 (N226, N1473);
	AND2X1 g_N1474 (N2233, N2582, N1474);
	AND2X1 g_N1475 (N157, N22, N1475);
	AND2X1 g_N1476 (N2898, N1862, N1476);
	BUFX2 g_N291 (N2018, N291);
	BUFX2 g_N1477 (N2592, N1477);
	BUFX2 g_N1478 (N1852, N1478);
	AND2X1 g_N1479 (N96, N213, N1479);
	BUFX2 g_N1480 (N1436, N1480);
	AND2X1 g_N1481 (N2872, N1730, N1481);
	INVX1 g_N1482 (N2491, N1482);
	INVX1 g_N1483 (N1047, N1483);
	INVX1 g_N1484 (N2940, N1484);
	BUFX2 g_N1485 (N2818, N1485);
	BUFX2 g_N1486 (N1159, N1486);
	BUFX2 g_N1487 (N2101, N1487);
	INVX1 g_N1488 (N3051, N1488);
	BUFX2 g_N292 (N689, N292);
	INVX1 g_N1489 (N2051, N1489);
	AND2X1 g_N1490 (N1496, N3387, N1490);
	BUFX2 g_N1491 (N1599, N1491);
	INVX1 g_N1492 (N1785, N1492);
	AND2X1 g_N1493 (N2778, N2736, N1493);
	INVX1 g_N1494 (N523, N1494);
	BUFX2 g_N1495 (N1651, N1495);
	INVX1 g_N1496 (N3403, N1496);
	AND2X1 g_N1497 (N713, N2415, N1497);
	AND2X1 g_N1498 (N665, N3418, N1498);
	INVX1 g_N1499 (N884, N1499);
	BUFX2 g_N1500 (N1788, N1500);
	AND2X1 g_N1501 (N418, N825, N1501);
	BUFX2 g_N1502 (N3067, N1502);
	INVX1 g_N1503 (N1086, N1503);
	INVX1 g_N1504 (N177, N1504);
	BUFX2 g_N1505 (N3883, N1505);
	AND2X1 g_N1506 (N726, N1753, N1506);
	AND2X1 g_N1507 (N1743, N2154, N1507);
	BUFX2 g_N293 (N1063, N293);
	INVX1 g_N1508 (N21, N1508);
	AND2X1 g_N1509 (N2830, N3095, N1509);
	BUFX2 g_N1510 (N2930, N1510);
	AND2X1 g_N1511 (N2926, N725, N1511);
	INVX1 g_N1512 (N3938, N1512);
	BUFX2 g_N1513 (N938, N1513);
	INVX1 g_N1514 (N1006, N1514);
	INVX1 g_N1515 (N3035, N1515);
	AND2X1 g_N1516 (N2738, N524, N1516);
	BUFX2 g_N1517 (N3919, N1517);
	AND2X1 g_N1518 (N2603, N2831, N1518);
	AND2X1 g_N1519 (N2276, N2264, N1519);
	INVX1 g_N1520 (N1252, N1520);
	INVX1 g_N1521 (N2700, N1521);
	BUFX2 g_N1522 (N2121, N1522);
	AND2X1 g_N1523 (N3798, N1460, N1523);
	BUFX2 g_N1524 (N2718, N1524);
	AND2X1 g_N1525 (N2724, N1561, N1525);
	BUFX2 g_N1526 (N1835, N1526);
	BUFX2 g_N1527 (N609, N1527);
	BUFX2 g_N1528 (N519, N1528);
	BUFX2 g_N1529 (N2610, N1529);
	INVX1 g_N1530 (N3015, N1530);
	INVX1 g_N1531 (N674, N1531);
	INVX1 g_N1532 (N2028, N1532);
	INVX1 g_N1533 (N58, N1533);
	INVX1 g_N1534 (N922, N1534);
	BUFX2 g_N1535 (N1095, N1535);
	INVX1 g_N1536 (N2404, N1536);
	AND2X1 g_N1537 (N1389, N2622, N1537);
	AND2X1 g_N1538 (N3846, N839, N1538);
	AND2X1 g_N1539 (N2136, N2971, N1539);
	BUFX2 g_N1540 (N1162, N1540);
	INVX1 g_N1541 (N2827, N1541);
	INVX1 g_N1542 (N2869, N1542);
	AND2X1 g_N1543 (N3640, N2571, N1543);
	INVX1 g_N1544 (N1416, N1544);
	INVX1 g_N1545 (N3672, N1545);
	INVX1 g_N1546 (N703, N1546);
	INVX1 g_N1547 (N3684, N1547);
	INVX1 g_N1548 (N1070, N1548);
	BUFX2 g_N1549 (N686, N1549);
	BUFX2 g_N1550 (N1455, N1550);
	BUFX2 g_N1551 (N2897, N1551);
	INVX1 g_N1552 (N2322, N1552);
	INVX1 g_N1553 (N1954, N1553);
	INVX1 g_N1554 (N3663, N1554);
	INVX1 g_N1555 (N2057, N1555);
	INVX1 g_N1556 (N5, N1556);
	INVX1 g_N1557 (N2661, N1557);
	INVX1 g_N1558 (N3192, N1558);
	AND2X1 g_N1559 (N2201, N1009, N1559);
	AND2X1 g_N1560 (N1619, N2133, N1560);
	INVX1 g_N1561 (N2528, N1561);
	INVX1 g_N1562 (N3619, N1562);
	AND2X1 g_N1563 (N1819, N3411, N1563);
	INVX1 g_N1564 (N3900, N1564);
	INVX1 g_N1565 (N1317, N1565);
	INVX1 g_N1566 (N1510, N1566);
	INVX1 g_N1567 (N2784, N1567);
	BUFX2 g_N1568 (N2962, N1568);
	INVX1 g_N1569 (N75, N1569);
	AND2X1 g_N1570 (N1764, N3427, N1570);
	INVX1 g_N1571 (N1375, N1571);
	BUFX2 g_N1572 (N3849, N1572);
	INVX1 g_N1573 (N146, N1573);
	INVX1 g_N1574 (N1272, N1574);
	BUFX2 g_N1575 (N1273, N1575);
	INVX1 g_N1576 (N2639, N1576);
	AND2X1 g_N1577 (N106, N117, N1577);
	BUFX2 g_N294 (N1946, N294);
	BUFX2 g_N1578 (N2917, N1578);
	INVX1 g_N1579 (N2400, N1579);
	AND2X1 g_N1580 (N3341, N1636, N1580);
	INVX1 g_N1581 (N117, N1581);
	AND2X1 g_N1582 (N2479, N575, N1582);
	INVX1 g_N1583 (N965, N1583);
	AND2X1 g_N1584 (N177, N188, N1584);
	INVX1 g_N1585 (N3258, N1585);
	INVX1 g_N1586 (N2475, N1586);
	AND2X1 g_N1587 (N2157, N1993, N1587);
	INVX1 g_N1588 (N2576, N1588);
	INVX1 g_N1589 (N462, N1589);
	BUFX2 g_N1590 (N3720, N1590);
	AND2X1 g_N1591 (N2485, N2494, N1591);
	BUFX2 g_N295 (N653, N295);
	BUFX2 g_N1592 (N1884, N1592);
	AND2X1 g_N1593 (N2053, N2033, N1593);
	AND2X1 g_N1594 (N2899, N3135, N1594);
	AND2X1 g_N1595 (N1130, N3251, N1595);
	INVX1 g_N1596 (N3561, N1596);
	BUFX2 g_N1597 (N800, N1597);
	INVX1 g_N1598 (N3225, N1598);
	AND2X1 g_N1599 (N105, N214, N1599);
	INVX1 g_N1600 (N232, N1600);
	INVX1 g_N1601 (N1082, N1601);
	BUFX2 g_N1602 (N2013, N1602);
	BUFX2 g_N1603 (N1886, N1603);
	AND2X1 g_N1604 (N3592, N2690, N1604);
	INVX1 g_N1605 (N49, N1605);
	INVX1 g_N1606 (N1761, N1606);
	BUFX2 g_N1607 (N1894, N1607);
	AND2X1 g_N1608 (N2403, N831, N1608);
	BUFX2 g_N296 (N2666, N296);
	INVX1 g_N1609 (N131, N1609);
	INVX1 g_N1610 (N1746, N1610);
	BUFX2 g_N1611 (N1837, N1611);
	AND2X1 g_N1612 (N1248, N755, N1612);
	INVX1 g_N1613 (N1923, N1613);
	INVX1 g_N1614 (N34, N1614);
	INVX1 g_N1615 (N462, N1615);
	BUFX2 g_N1616 (N3203, N1616);
	INVX1 g_N1617 (N3558, N1617);
	AND2X1 g_N1618 (N3693, N1548, N1618);
	INVX1 g_N1619 (N3252, N1619);
	INVX1 g_N1620 (N2927, N1620);
	BUFX2 g_N297 (N1989, N297);
	BUFX2 g_N1621 (N2118, N1621);
	BUFX2 g_N1622 (N2546, N1622);
	INVX1 g_N1623 (N2810, N1623);
	AND2X1 g_N1624 (N607, N450, N1624);
	INVX1 g_N1625 (N142, N1625);
	AND2X1 g_N1626 (N2554, N3249, N1626);
	BUFX2 g_N298 (N2037, N298);
	INVX1 g_N1627 (N2432, N1627);
	BUFX2 g_N1628 (N3375, N1628);
	INVX1 g_N1629 (N85, N1629);
	AND2X1 g_N1630 (N3351, N3676, N1630);
	AND2X1 g_N1631 (N2454, N3476, N1631);
	INVX1 g_N1632 (N2002, N1632);
	BUFX2 g_N1633 (N754, N1633);
	INVX1 g_N1634 (N645, N1634);
	AND2X1 g_N1635 (N589, N3734, N1635);
	INVX1 g_N1636 (N1778, N1636);
	INVX1 g_N1637 (N2430, N1637);
	INVX1 g_N1638 (N1057, N1638);
	INVX1 g_N1639 (N2487, N1639);
	AND2X1 g_N1640 (N3913, N2862, N1640);
	INVX1 g_N1641 (N541, N1641);
	INVX1 g_N1642 (N1858, N1642);
	INVX1 g_N1643 (N1302, N1643);
	AND2X1 g_N1644 (N3483, N1746, N1644);
	BUFX2 g_N1645 (N3076, N1645);
	AND2X1 g_N1646 (N225, N87, N1646);
	BUFX2 g_N1647 (N2480, N1647);
	AND2X1 g_N1648 (N2819, N434, N1648);
	INVX1 g_N1649 (N1467, N1649);
	AND2X1 g_N1650 (N1699, N3144, N1650);
	AND2X1 g_N1651 (N3373, N806, N1651);
	AND2X1 g_N1652 (N926, N3549, N1652);
	BUFX2 g_N1653 (N2271, N1653);
	AND2X1 g_N1654 (N68, N160, N1654);
	AND2X1 g_N1655 (N2169, N1008, N1655);
	INVX1 g_N1656 (N3094, N1656);
	INVX1 g_N1657 (N1868, N1657);
	AND2X1 g_N1658 (N3090, N3484, N1658);
	INVX1 g_N1659 (N2309, N1659);
	BUFX2 g_N1660 (N3642, N1660);
	AND2X1 g_N1661 (N3571, N1710, N1661);
	BUFX2 g_N1662 (N1387, N1662);
	INVX1 g_N1663 (N1045, N1663);
	AND2X1 g_N1664 (N3112, N720, N1664);
	AND2X1 g_N1665 (N1974, N1188, N1665);
	AND2X1 g_N1666 (N2585, N1155, N1666);
	INVX1 g_N1667 (N3200, N1667);
	INVX1 g_N1668 (N930, N1668);
	AND2X1 g_N1669 (N1572, N2498, N1669);
	INVX1 g_N1670 (N2021, N1670);
	INVX1 g_N1671 (N1602, N1671);
	INVX1 g_N1672 (N2182, N1672);
	AND2X1 g_N1673 (N2573, N3103, N1673);
	BUFX2 g_N1674 (N2341, N1674);
	AND2X1 g_N1675 (N1562, N2638, N1675);
	INVX1 g_N1676 (N1945, N1676);
	INVX1 g_N1677 (N2473, N1677);
	AND2X1 g_N1678 (N2005, N829, N1678);
	AND2X1 g_N1679 (N2425, N765, N1679);
	AND2X1 g_N1680 (N3013, N2426, N1680);
	BUFX2 g_N1681 (N3189, N1681);
	BUFX2 g_N1682 (N2943, N1682);
	BUFX2 g_N1683 (N1359, N1683);
	BUFX2 g_N1684 (N1994, N1684);
	AND2X1 g_N1685 (N1547, N3694, N1685);
	AND2X1 g_N1686 (N1271, N1824, N1686);
	INVX1 g_N1687 (N945, N1687);
	AND2X1 g_N1688 (N245, N8, N1688);
	INVX1 g_N1689 (N3656, N1689);
	AND2X1 g_N1690 (N3853, N2725, N1690);
	BUFX2 g_N1691 (N635, N1691);
	INVX1 g_N1692 (N236, N1692);
	INVX1 g_N1693 (N717, N1693);
	INVX1 g_N1694 (N13, N1694);
	AND2X1 g_N1695 (N2865, N1880, N1695);
	AND2X1 g_N1696 (N2944, N2702, N1696);
	BUFX2 g_N1697 (N2530, N1697);
	BUFX2 g_N1698 (N1820, N1698);
	BUFX2 g_N1699 (N1316, N1699);
	INVX1 g_N1700 (N615, N1700);
	AND2X1 g_N1701 (N763, N565, N1701);
	AND2X1 g_N1702 (N3134, N423, N1702);
	INVX1 g_N1703 (N2684, N1703);
	BUFX2 g_N299 (N821, N299);
	BUFX2 g_N1704 (N2617, N1704);
	AND2X1 g_N1705 (N995, N1154, N1705);
	INVX1 g_N1706 (N3631, N1706);
	INVX1 g_N1707 (N3389, N1707);
	BUFX2 g_N300 (N2651, N300);
	INVX1 g_N1708 (N2024, N1708);
	BUFX2 g_N1709 (N2164, N1709);
	INVX1 g_N1710 (N169, N1710);
	INVX1 g_N1711 (N2282, N1711);
	INVX1 g_N1712 (N1200, N1712);
	INVX1 g_N1713 (N88, N1713);
	AND2X1 g_N1714 (N1196, N182, N1714);
	AND2X1 g_N1715 (N2110, N3681, N1715);
	AND2X1 g_N1716 (N1898, N1900, N1716);
	BUFX2 g_N1717 (N1309, N1717);
	INVX1 g_N1718 (N1007, N1718);
	AND2X1 g_N1719 (N195, N181, N1719);
	BUFX2 g_N301 (N1449, N301);
	INVX1 g_N1720 (N3933, N1720);
	INVX1 g_N1721 (N72, N1721);
	AND2X1 g_N1722 (N253, N36, N1722);
	AND2X1 g_N1723 (N1003, N1356, N1723);
	AND2X1 g_N1724 (N3861, N2834, N1724);
	INVX1 g_N1725 (N3018, N1725);
	INVX1 g_N1726 (N3422, N1726);
	AND2X1 g_N1727 (N1199, N2757, N1727);
	AND2X1 g_N1728 (N3678, N956, N1728);
	BUFX2 g_N1729 (N3741, N1729);
	INVX1 g_N1730 (N16, N1730);
	INVX1 g_N1731 (N941, N1731);
	INVX1 g_N1732 (N2350, N1732);
	INVX1 g_N1733 (N1265, N1733);
	INVX1 g_N1734 (N503, N1734);
	AND2X1 g_N1735 (N85, N42, N1735);
	INVX1 g_N1736 (N2456, N1736);
	AND2X1 g_N1737 (N208, N176, N1737);
	INVX1 g_N1738 (N159, N1738);
	AND2X1 g_N1739 (N1285, N3314, N1739);
	INVX1 g_N1740 (N3549, N1740);
	INVX1 g_N1741 (N2895, N1741);
	BUFX2 g_N1742 (N2127, N1742);
	INVX1 g_N1743 (N972, N1743);
	BUFX2 g_N1744 (N962, N1744);
	INVX1 g_N1745 (N1358, N1745);
	BUFX2 g_N1746 (N1675, N1746);
	INVX1 g_N1747 (N2306, N1747);
	BUFX2 g_N1748 (N1580, N1748);
	AND2X1 g_N1749 (N3844, N1495, N1749);
	AND2X1 g_N1750 (N1576, N2224, N1750);
	BUFX2 g_N1751 (N1461, N1751);
	INVX1 g_N1752 (N796, N1752);
	INVX1 g_N1753 (N3535, N1753);
	INVX1 g_N1754 (N2899, N1754);
	BUFX2 g_N1755 (N2499, N1755);
	INVX1 g_N1756 (N835, N1756);
	AND2X1 g_N1757 (N3688, N2985, N1757);
	AND2X1 g_N1758 (N2611, N1589, N1758);
	BUFX2 g_N1759 (N3702, N1759);
	INVX1 g_N1760 (N2416, N1760);
	BUFX2 g_N1761 (N2113, N1761);
	INVX1 g_N1762 (N2730, N1762);
	BUFX2 g_N1763 (N399, N1763);
	INVX1 g_N1764 (N798, N1764);
	BUFX2 g_N302 (N657, N302);
	BUFX2 g_N1765 (N1511, N1765);
	INVX1 g_N1766 (N112, N1766);
	AND2X1 g_N1767 (N2317, N2392, N1767);
	INVX1 g_N1768 (N1477, N1768);
	INVX1 g_N1769 (N3142, N1769);
	BUFX2 g_N1770 (N1065, N1770);
	INVX1 g_N1771 (N1144, N1771);
	BUFX2 g_N1772 (N1493, N1772);
	INVX1 g_N1773 (N3613, N1773);
	INVX1 g_N1774 (N242, N1774);
	AND2X1 g_N1775 (N778, N1211, N1775);
	AND2X1 g_N1776 (N1337, N2046, N1776);
	BUFX2 g_N1777 (N1004, N1777);
	BUFX2 g_N1778 (N3796, N1778);
	INVX1 g_N1779 (N1326, N1779);
	AND2X1 g_N1780 (N873, N1713, N1780);
	INVX1 g_N1781 (N3549, N1781);
	INVX1 g_N1782 (N642, N1782);
	AND2X1 g_N1783 (N1331, N1792, N1783);
	INVX1 g_N1784 (N221, N1784);
	BUFX2 g_N1785 (N714, N1785);
	INVX1 g_N1786 (N690, N1786);
	BUFX2 g_N1787 (N2001, N1787);
	AND2X1 g_N1788 (N843, N1821, N1788);
	INVX1 g_N1789 (N134, N1789);
	BUFX2 g_N1790 (N2234, N1790);
	INVX1 g_N1791 (N2967, N1791);
	INVX1 g_N1792 (N2293, N1792);
	INVX1 g_N1793 (N2285, N1793);
	INVX1 g_N1794 (N224, N1794);
	AND2X1 g_N1795 (N865, N3622, N1795);
	AND2X1 g_N1796 (N3323, N1092, N1796);
	INVX1 g_N1797 (N82, N1797);
	INVX1 g_N1798 (N3840, N1798);
	AND2X1 g_N1799 (N1598, N3889, N1799);
	BUFX2 g_N1800 (N2629, N1800);
	INVX1 g_N1801 (N1831, N1801);
	BUFX2 g_N1802 (N2608, N1802);
	INVX1 g_N1803 (N1988, N1803);
	AND2X1 g_N1804 (N3823, N2817, N1804);
	INVX1 g_N1805 (N2870, N1805);
	BUFX2 g_N303 (N3723, N303);
	BUFX2 g_N1806 (N2768, N1806);
	AND2X1 g_N1807 (N2213, N1238, N1807);
	AND2X1 g_N1808 (N1304, N629, N1808);
	BUFX2 g_N1809 (N2279, N1809);
	AND2X1 g_N1810 (N2956, N3450, N1810);
	BUFX2 g_N304 (N3532, N304);
	BUFX2 g_N1811 (N3297, N1811);
	INVX1 g_N1812 (N500, N1812);
	BUFX2 g_N1813 (N612, N1813);
	AND2X1 g_N1814 (N769, N992, N1814);
	INVX1 g_N1815 (N1653, N1815);
	AND2X1 g_N1816 (N1960, N1375, N1816);
	INVX1 g_N1817 (N154, N1817);
	AND2X1 g_N1818 (N1392, N2261, N1818);
	BUFX2 g_N1819 (N780, N1819);
	AND2X1 g_N1820 (N1520, N718, N1820);
	INVX1 g_N1821 (N1487, N1821);
	INVX1 g_N1822 (N572, N1822);
	AND2X1 g_N1823 (N419, N2484, N1823);
	INVX1 g_N1824 (N1338, N1824);
	INVX1 g_N1825 (N1055, N1825);
	BUFX2 g_N1826 (N1215, N1826);
	INVX1 g_N1827 (N2208, N1827);
	INVX1 g_N1828 (N622, N1828);
	INVX1 g_N1829 (N703, N1829);
	BUFX2 g_N1830 (N1807, N1830);
	BUFX2 g_N1831 (N3813, N1831);
	BUFX2 g_N1832 (N3091, N1832);
	AND2X1 g_N1833 (N1431, N1334, N1833);
	INVX1 g_N1834 (N2134, N1834);
	AND2X1 g_N1835 (N2041, N1144, N1835);
	BUFX2 g_N305 (N1257, N305);
	AND2X1 g_N1836 (N1043, N3479, N1836);
	BUFX2 g_N306 (N1134, N306);
	AND2X1 g_N1837 (N2267, N2347, N1837);
	BUFX2 g_N1838 (N2191, N1838);
	AND2X1 g_N1839 (N2634, N2774, N1839);
	INVX1 g_N1840 (N2933, N1840);
	AND2X1 g_N1841 (N1275, N1922, N1841);
	BUFX2 g_N1842 (N1618, N1842);
	AND2X1 g_N1843 (N2500, N3151, N1843);
	INVX1 g_N1844 (N2492, N1844);
	AND2X1 g_N1845 (N2873, N944, N1845);
	AND2X1 g_N1846 (N10, N112, N1846);
	INVX1 g_N1847 (N2614, N1847);
	AND2X1 g_N1848 (N3842, N679, N1848);
	BUFX2 g_N1849 (N974, N1849);
	INVX1 g_N1850 (N3548, N1850);
	INVX1 g_N1851 (N1452, N1851);
	AND2X1 g_N1852 (N479, N3851, N1852);
	AND2X1 g_N1853 (N2856, N3258, N1853);
	INVX1 g_N1854 (N847, N1854);
	INVX1 g_N1855 (N3036, N1855);
	INVX1 g_N1856 (N1023, N1856);
	AND2X1 g_N1857 (N2329, N1094, N1857);
	BUFX2 g_N1858 (N1361, N1858);
	INVX1 g_N1859 (N3884, N1859);
	AND2X1 g_N1860 (N3128, N1662, N1860);
	BUFX2 g_N1861 (N3574, N1861);
	BUFX2 g_N1862 (N2959, N1862);
	BUFX2 g_N1863 (N3021, N1863);
	INVX1 g_N1864 (N176, N1864);
	AND2X1 g_N1865 (N2286, N529, N1865);
	INVX1 g_N1866 (N2406, N1866);
	BUFX2 g_N1867 (N3461, N1867);
	BUFX2 g_N1868 (N1234, N1868);
	INVX1 g_N1869 (N1431, N1869);
	AND2X1 g_N1870 (N2543, N3442, N1870);
	BUFX2 g_N1871 (N661, N1871);
	BUFX2 g_N1872 (N1380, N1872);
	BUFX2 g_N1873 (N1443, N1873);
	AND2X1 g_N1874 (N2103, N1607, N1874);
	INVX1 g_N1875 (N1241, N1875);
	INVX1 g_N1876 (N1495, N1876);
	BUFX2 g_N1877 (N1665, N1877);
	BUFX2 g_N1878 (N676, N1878);
	BUFX2 g_N307 (N662, N307);
	INVX1 g_N1879 (N1933, N1879);
	BUFX2 g_N1880 (N1679, N1880);
	INVX1 g_N1881 (N111, N1881);
	INVX1 g_N1882 (N1452, N1882);
	INVX1 g_N1883 (N738, N1883);
	AND2X1 g_N1884 (N35, N40, N1884);
	AND2X1 g_N1885 (N2092, N3625, N1885);
	AND2X1 g_N1886 (N2949, N1542, N1886);
	AND2X1 g_N1887 (N1971, N692, N1887);
	AND2X1 g_N1888 (N1861, N1771, N1888);
	INVX1 g_N1889 (N2754, N1889);
	INVX1 g_N1890 (N1074, N1890);
	AND2X1 g_N1891 (N2023, N3023, N1891);
	INVX1 g_N1892 (N457, N1892);
	INVX1 g_N1893 (N31, N1893);
	AND2X1 g_N1894 (N2062, N2167, N1894);
	BUFX2 g_N1895 (N2372, N1895);
	INVX1 g_N1896 (N3619, N1896);
	INVX1 g_N1897 (N1329, N1897);
	INVX1 g_N1898 (N3343, N1898);
	BUFX2 g_N1899 (N1197, N1899);
	INVX1 g_N1900 (N1409, N1900);
	AND2X1 g_N1901 (N3041, N3099, N1901);
	BUFX2 g_N1902 (N999, N1902);
	BUFX2 g_N1903 (N3929, N1903);
	INVX1 g_N1904 (N1252, N1904);
	BUFX2 g_N1905 (N2682, N1905);
	BUFX2 g_N1906 (N986, N1906);
	AND2X1 g_N1907 (N616, N2273, N1907);
	INVX1 g_N1908 (N2385, N1908);
	INVX1 g_N1909 (N1167, N1909);
	INVX1 g_N1910 (N1044, N1910);
	INVX1 g_N1911 (N2606, N1911);
	AND2X1 g_N1912 (N2497, N2155, N1912);
	BUFX2 g_N1913 (N2979, N1913);
	BUFX2 g_N1914 (N2513, N1914);
	INVX1 g_N1915 (N1062, N1915);
	INVX1 g_N1916 (N1930, N1916);
	AND2X1 g_N1917 (N3198, N1530, N1917);
	AND2X1 g_N1918 (N2545, N1873, N1918);
	INVX1 g_N1919 (N618, N1919);
	BUFX2 g_N1920 (N710, N1920);
	INVX1 g_N1921 (N129, N1921);
	INVX1 g_N1922 (N1505, N1922);
	BUFX2 g_N1923 (N561, N1923);
	AND2X1 g_N1924 (N1997, N1798, N1924);
	BUFX2 g_N1925 (N1696, N1925);
	BUFX2 g_N1926 (N2871, N1926);
	INVX1 g_N1927 (N3402, N1927);
	AND2X1 g_N1928 (N3374, N2068, N1928);
	AND2X1 g_N1929 (N934, N3465, N1929);
	BUFX2 g_N1930 (N604, N1930);
	INVX1 g_N1931 (N2465, N1931);
	AND2X1 g_N1932 (N1762, N1950, N1932);
	BUFX2 g_N1933 (N3925, N1933);
	AND2X1 g_N1934 (N1364, N474, N1934);
	INVX1 g_N1935 (N2154, N1935);
	AND2X1 g_N1936 (N1681, N3029, N1936);
	AND2X1 g_N1937 (N2093, N2371, N1937);
	AND2X1 g_N1938 (N2241, N552, N1938);
	AND2X1 g_N1939 (N3878, N2595, N1939);
	AND2X1 g_N1940 (N2581, N2887, N1940);
	AND2X1 g_N1941 (N1421, N1784, N1941);
	AND2X1 g_N1942 (N3597, N3012, N1942);
	INVX1 g_N1943 (N1178, N1943);
	BUFX2 g_N1944 (N2448, N1944);
	BUFX2 g_N1945 (N3825, N1945);
	BUFX2 g_N1946 (N1138, N1946);
	INVX1 g_N1947 (N2684, N1947);
	INVX1 g_N1948 (N2160, N1948);
	INVX1 g_N1949 (N2050, N1949);
	BUFX2 g_N308 (N2123, N308);
	INVX1 g_N1950 (N3207, N1950);
	AND2X1 g_N1951 (N3139, N1169, N1951);
	AND2X1 g_N1952 (N205, N228, N1952);
	INVX1 g_N1953 (N35, N1953);
	BUFX2 g_N1954 (N3460, N1954);
	BUFX2 g_N1955 (N1924, N1955);
	INVX1 g_N1956 (N4, N1956);
	BUFX2 g_N1957 (N2367, N1957);
	BUFX2 g_N1958 (N1932, N1958);
	BUFX2 g_N309 (N2707, N309);
	INVX1 g_N1959 (N113, N1959);
	INVX1 g_N1960 (N3410, N1960);
	AND2X1 g_N1961 (N1615, N1979, N1961);
	INVX1 g_N1962 (N1404, N1962);
	INVX1 g_N1963 (N229, N1963);
	BUFX2 g_N1964 (N2993, N1964);
	BUFX2 g_N1965 (N1595, N1965);
	INVX1 g_N1966 (N1495, N1966);
	BUFX2 g_N1967 (N1507, N1967);
	BUFX2 g_N1968 (N2031, N1968);
	AND2X1 g_N1969 (N2635, N3222, N1969);
	INVX1 g_N1970 (N3710, N1970);
	INVX1 g_N1971 (N150, N1971);
	INVX1 g_N1972 (N218, N1972);
	INVX1 g_N1973 (N546, N1973);
	INVX1 g_N1974 (N1057, N1974);
	BUFX2 g_N1975 (N2821, N1975);
	INVX1 g_N1976 (N71, N1976);
	INVX1 g_N1977 (N739, N1977);
	AND2X1 g_N1978 (N3696, N2134, N1978);
	INVX1 g_N1979 (N3082, N1979);
	BUFX2 g_N1980 (N853, N1980);
	AND2X1 g_N1981 (N159, N141, N1981);
	BUFX2 g_N1982 (N3482, N1982);
	BUFX2 g_N1983 (N3263, N1983);
	INVX1 g_N1984 (N1027, N1984);
	AND2X1 g_N1985 (N227, N65, N1985);
	BUFX2 g_N1986 (N2883, N1986);
	INVX1 g_N1987 (N1681, N1987);
	BUFX2 g_N1988 (N3726, N1988);
	BUFX2 g_N1989 (N1685, N1989);
	INVX1 g_N1990 (N501, N1990);
	BUFX2 g_N1991 (N3079, N1991);
	BUFX2 g_N1992 (N3448, N1992);
	INVX1 g_N1993 (N437, N1993);
	AND2X1 g_N1994 (N6, N53, N1994);
	INVX1 g_N1995 (N961, N1995);
	BUFX2 g_N1996 (N3765, N1996);
	INVX1 g_N1997 (N1878, N1997);
	BUFX2 g_N310 (N2345, N310);
	INVX1 g_N1998 (N3433, N1998);
	INVX1 g_N1999 (N1647, N1999);
	INVX1 g_N2000 (N3238, N2000);
	AND2X1 g_N2001 (N3620, N2884, N2001);
	BUFX2 g_N2002 (N1243, N2002);
	AND2X1 g_N2003 (N3492, N3945, N2003);
	INVX1 g_N2004 (N220, N2004);
	INVX1 g_N2005 (N1965, N2005);
	AND2X1 g_N2006 (N201, N49, N2006);
	BUFX2 g_N2007 (N2589, N2007);
	BUFX2 g_N2008 (N3240, N2008);
	INVX1 g_N2009 (N3573, N2009);
	AND2X1 g_N2010 (N2553, N3347, N2010);
	AND2X1 g_N2011 (N3037, N1179, N2011);
	AND2X1 g_N2012 (N3345, N2940, N2012);
	AND2X1 g_N2013 (N62, N132, N2013);
	AND2X1 g_N2014 (N1500, N3202, N2014);
	INVX1 g_N2015 (N1755, N2015);
	BUFX2 g_N311 (N1551, N311);
	AND2X1 g_N2016 (N3607, N1477, N2016);
	INVX1 g_N2017 (N1090, N2017);
	BUFX2 g_N2018 (N3342, N2018);
	BUFX2 g_N2019 (N2360, N2019);
	BUFX2 g_N2020 (N2712, N2020);
	BUFX2 g_N2021 (N1678, N2021);
	BUFX2 g_N312 (N3453, N312);
	INVX1 g_N2022 (N155, N2022);
	INVX1 g_N2023 (N103, N2023);
	BUFX2 g_N2024 (N1885, N2024);
	INVX1 g_N2025 (N3629, N2025);
	INVX1 g_N2026 (N3051, N2026);
	AND2X1 g_N2027 (N1889, N2769, N2027);
	BUFX2 g_N2028 (N3701, N2028);
	AND2X1 g_N2029 (N2852, N849, N2029);
	BUFX2 g_N313 (N3268, N313);
	INVX1 g_N2030 (N2061, N2030);
	AND2X1 g_N2031 (N3885, N1752, N2031);
	BUFX2 g_N2032 (N1156, N2032);
	INVX1 g_N2033 (N3673, N2033);
	INVX1 g_N2034 (N3217, N2034);
	BUFX2 g_N2035 (N2727, N2035);
	INVX1 g_N2036 (N3714, N2036);
	BUFX2 g_N2037 (N2823, N2037);
	BUFX2 g_N2038 (N3655, N2038);
	AND2X1 g_N2039 (N1093, N3477, N2039);
	INVX1 g_N2040 (N76, N2040);
	BUFX2 g_N314 (N559, N314);
	INVX1 g_N2041 (N1861, N2041);
	INVX1 g_N2042 (N1081, N2042);
	INVX1 g_N2043 (N654, N2043);
	INVX1 g_N2044 (N1529, N2044);
	BUFX2 g_N2045 (N2106, N2045);
	INVX1 g_N2046 (N1578, N2046);
	AND2X1 g_N2047 (N3116, N1671, N2047);
	INVX1 g_N2048 (N409, N2048);
	BUFX2 g_N2049 (N1297, N2049);
	BUFX2 g_N2050 (N1231, N2050);
	BUFX2 g_N2051 (N1434, N2051);
	AND2X1 g_N2052 (N2808, N2211, N2052);
	INVX1 g_N2053 (N3903, N2053);
	AND2X1 g_N2054 (N2204, N2941, N2054);
	INVX1 g_N2055 (N2561, N2055);
	INVX1 g_N2056 (N540, N2056);
	BUFX2 g_N2057 (N3206, N2057);
	INVX1 g_N2058 (N3867, N2058);
	INVX1 g_N2059 (N1903, N2059);
	BUFX2 g_N315 (N711, N315);
	INVX1 g_N2060 (N3386, N2060);
	BUFX2 g_N2061 (N2115, N2061);
	INVX1 g_N2062 (N2714, N2062);
	AND2X1 g_N2063 (N748, N3177, N2063);
	INVX1 g_N2064 (N15, N2064);
	BUFX2 g_N2065 (N2988, N2065);
	INVX1 g_N2066 (N2785, N2066);
	BUFX2 g_N2067 (N2825, N2067);
	INVX1 g_N2068 (N2740, N2068);
	INVX1 g_N2069 (N1385, N2069);
	AND2X1 g_N2070 (N2058, N3616, N2070);
	BUFX2 g_N316 (N3528, N316);
	BUFX2 g_N2071 (N826, N2071);
	INVX1 g_N2072 (N1872, N2072);
	AND2X1 g_N2073 (N2809, N693, N2073);
	INVX1 g_N2074 (N106, N2074);
	INVX1 g_N2075 (N1607, N2075);
	INVX1 g_N2076 (N243, N2076);
	AND2X1 g_N2077 (N44, N83, N2077);
	BUFX2 g_N2078 (N2532, N2078);
	INVX1 g_N2079 (N3258, N2079);
	BUFX2 g_N2080 (N1068, N2080);
	OR2X1 g_N2081 (N2540, N2183, N2081);
	AND2X1 g_N2082 (N3542, N2146, N2082);
	INVX1 g_N2083 (N1310, N2083);
	INVX1 g_N2084 (N3420, N2084);
	INVX1 g_N2085 (N3615, N2085);
	INVX1 g_N2086 (N1071, N2086);
	INVX1 g_N2087 (N1335, N2087);
	BUFX2 g_N2088 (N3289, N2088);
	INVX1 g_N2089 (N70, N2089);
	INVX1 g_N2090 (N389, N2090);
	INVX1 g_N2091 (N90, N2091);
	INVX1 g_N2092 (N25, N2092);
	INVX1 g_N2093 (N2895, N2093);
	INVX1 g_N2094 (N2627, N2094);
	AND2X1 g_N2095 (N1801, N1822, N2095);
	AND2X1 g_N2096 (N797, N808, N2096);
	BUFX2 g_N2097 (N3766, N2097);
	BUFX2 g_N2098 (N2359, N2098);
	INVX1 g_N2099 (N3088, N2099);
	BUFX2 g_N2100 (N2082, N2100);
	AND2X1 g_N2101 (N242, N80, N2101);
	AND2X1 g_N2102 (N2205, N601, N2102);
	INVX1 g_N2103 (N2519, N2103);
	INVX1 g_N2104 (N1996, N2104);
	BUFX2 g_N2105 (N861, N2105);
	AND2X1 g_N2106 (N1191, N1774, N2106);
	INVX1 g_N2107 (N1067, N2107);
	INVX1 g_N2108 (N2981, N2108);
	BUFX2 g_N2109 (N660, N2109);
	INVX1 g_N2110 (N3463, N2110);
	INVX1 g_N2111 (N963, N2111);
	INVX1 g_N2112 (N976, N2112);
	AND2X1 g_N2113 (N3359, N3859, N2113);
	AND2X1 g_N2114 (N3309, N1999, N2114);
	AND2X1 g_N2115 (N2923, N697, N2115);
	INVX1 g_N2116 (N3288, N2116);
	INVX1 g_N2117 (N3332, N2117);
	AND2X1 g_N2118 (N1015, N3553, N2118);
	INVX1 g_N2119 (N1168, N2119);
	INVX1 g_N2120 (N2293, N2120);
	AND2X1 g_N2121 (N2129, N2409, N2121);
	INVX1 g_N2122 (N2531, N2122);
	BUFX2 g_N2123 (N1501, N2123);
	INVX1 g_N2124 (N3311, N2124);
	AND2X1 g_N2125 (N1250, N1906, N2125);
	AND2X1 g_N2126 (N1006, N3863, N2126);
	AND2X1 g_N2127 (N12, N7, N2127);
	AND2X1 g_N2128 (N3174, N2547, N2128);
	INVX1 g_N2129 (N1048, N2129);
	AND2X1 g_N2130 (N2746, N517, N2130);
	BUFX2 g_N2131 (N2495, N2131);
	AND2X1 g_N2132 (N95, N210, N2132);
	INVX1 g_N2133 (N927, N2133);
	BUFX2 g_N2134 (N3467, N2134);
	BUFX2 g_N2135 (N2466, N2135);
	INVX1 g_N2136 (N3767, N2136);
	BUFX2 g_N2137 (N417, N2137);
	BUFX2 g_N2138 (N2014, N2138);
	AND2X1 g_N2139 (N5, N60, N2139);
	BUFX2 g_N2140 (N3178, N2140);
	INVX1 g_N2141 (N1074, N2141);
	BUFX2 g_N2142 (N2326, N2142);
	AND2X1 g_N2143 (N1471, N1433, N2143);
	BUFX2 g_N2144 (N698, N2144);
	AND2X1 g_N2145 (N3415, N683, N2145);
	BUFX2 g_N2146 (N1151, N2146);
	AND2X1 g_N2147 (N2695, N792, N2147);
	AND2X1 g_N2148 (N1378, N3421, N2148);
	BUFX2 g_N2149 (N3318, N2149);
	AND2X1 g_N2150 (N3214, N864, N2150);
	AND2X1 g_N2151 (N3280, N403, N2151);
	BUFX2 g_N2152 (N2340, N2152);
	BUFX2 g_N2153 (N3401, N2153);
	BUFX2 g_N2154 (N2516, N2154);
	INVX1 g_N2155 (N2146, N2155);
	BUFX2 g_N2156 (N3804, N2156);
	INVX1 g_N2157 (N922, N2157);
	BUFX2 g_N2158 (N1414, N2158);
	INVX1 g_N2159 (N2671, N2159);
	BUFX2 g_N2160 (N1135, N2160);
	AND2X1 g_N2161 (N2583, N2247, N2161);
	BUFX2 g_N2162 (N2782, N2162);
	AND2X1 g_N2163 (N2854, N1641, N2163);
	AND2X1 g_N2164 (N411, N3488, N2164);
	BUFX2 g_N2165 (N3106, N2165);
	INVX1 g_N2166 (N1568, N2166);
	INVX1 g_N2167 (N2627, N2167);
	AND2X1 g_N2168 (N1581, N2074, N2168);
	INVX1 g_N2169 (N2071, N2169);
	BUFX2 g_N2170 (N2504, N2170);
	INVX1 g_N2171 (N1407, N2171);
	BUFX2 g_N2172 (N1587, N2172);
	AND2X1 g_N2173 (N2444, N1102, N2173);
	INVX1 g_N2174 (N450, N2174);
	INVX1 g_N2175 (N1312, N2175);
	INVX1 g_N2176 (N1480, N2176);
	INVX1 g_N2177 (N1395, N2177);
	INVX1 g_N2178 (N1107, N2178);
	INVX1 g_N2179 (N751, N2179);
	INVX1 g_N2180 (N1991, N2180);
	BUFX2 g_N2181 (N2578, N2181);
	BUFX2 g_N2182 (N3781, N2182);
	BUFX2 g_N317 (N3165, N317);
	BUFX2 g_N2183 (N3243, N2183);
	INVX1 g_N2184 (N659, N2184);
	AND2X1 g_N2185 (N1725, N2909, N2185);
	BUFX2 g_N2186 (N3539, N2186);
	BUFX2 g_N2187 (N761, N2187);
	AND2X1 g_N2188 (N1310, N2637, N2188);
	INVX1 g_N2189 (N3080, N2189);
	AND2X1 g_N2190 (N184, N229, N2190);
	AND2X1 g_N2191 (N2674, N1294, N2191);
	AND2X1 g_N2192 (N3719, N1545, N2192);
	INVX1 g_N2193 (N967, N2193);
	INVX1 g_N2194 (N122, N2194);
	BUFX2 g_N2195 (N2820, N2195);
	BUFX2 g_N2196 (N3526, N2196);
	AND2X1 g_N2197 (N3262, N702, N2197);
	BUFX2 g_N2198 (N951, N2198);
	INVX1 g_N2199 (N2487, N2199);
	BUFX2 g_N2200 (N3506, N2200);
	INVX1 g_N2201 (N820, N2201);
	AND2X1 g_N2202 (N1018, N1766, N2202);
	BUFX2 g_N2203 (N1981, N2203);
	INVX1 g_N2204 (N912, N2204);
	INVX1 g_N2205 (N637, N2205);
	INVX1 g_N2206 (N1241, N2206);
	BUFX2 g_N2207 (N2126, N2207);
	BUFX2 g_N2208 (N1426, N2208);
	BUFX2 g_N2209 (N1325, N2209);
	INVX1 g_N2210 (N2748, N2210);
	INVX1 g_N2211 (N3663, N2211);
	BUFX2 g_N318 (N663, N318);
	BUFX2 g_N2212 (N2538, N2212);
	INVX1 g_N2213 (N119, N2213);
	INVX1 g_N2214 (N1039, N2214);
	BUFX2 g_N2215 (N1630, N2215);
	BUFX2 g_N2216 (N1276, N2216);
	BUFX2 g_N2217 (N2482, N2217);
	BUFX2 g_N319 (N3237, N319);
	INVX1 g_N2218 (N838, N2218);
	INVX1 g_N2219 (N499, N2219);
	INVX1 g_N2220 (N3887, N2220);
	AND2X1 g_N2221 (N1569, N2536, N2221);
	INVX1 g_N2222 (N699, N2222);
	AND2X1 g_N2223 (N113, N23, N2223);
	BUFX2 g_N2224 (N3869, N2224);
	INVX1 g_N2225 (N27, N2225);
	INVX1 g_N2226 (N3336, N2226);
	AND2X1 g_N2227 (N998, N1362, N2227);
	AND2X1 g_N2228 (N893, N2890, N2228);
	AND2X1 g_N2229 (N52, N233, N2229);
	INVX1 g_N2230 (N2699, N2230);
	AND2X1 g_N2231 (N3060, N1470, N2231);
	BUFX2 g_N2232 (N712, N2232);
	INVX1 g_N2233 (N3576, N2233);
	AND2X1 g_N2234 (N2751, N2681, N2234);
	INVX1 g_N2235 (N2743, N2235);
	BUFX2 g_N2236 (N1122, N2236);
	AND2X1 g_N2237 (N547, N2009, N2237);
	AND2X1 g_N2238 (N1972, N2396, N2238);
	AND2X1 g_N2239 (N2572, N2319, N2239);
	BUFX2 g_N2240 (N2620, N2240);
	BUFX2 g_N320 (N2098, N320);
	BUFX2 g_N2241 (N1796, N2241);
	INVX1 g_N2242 (N3641, N2242);
	INVX1 g_N2243 (N3548, N2243);
	INVX1 g_N2244 (N245, N2244);
	AND2X1 g_N2245 (N164, N25, N2245);
	INVX1 g_N2246 (N2394, N2246);
	INVX1 g_N2247 (N2960, N2247);
	BUFX2 g_N2248 (N2389, N2248);
	BUFX2 g_N2249 (N1139, N2249);
	INVX1 g_N2250 (N120, N2250);
	BUFX2 g_N2251 (N388, N2251);
	INVX1 g_N2252 (N2381, N2252);
	INVX1 g_N2253 (N2827, N2253);
	INVX1 g_N2254 (N2758, N2254);
	INVX1 g_N2255 (N195, N2255);
	INVX1 g_N2256 (N941, N2256);
	BUFX2 g_N2257 (N1750, N2257);
	BUFX2 g_N2258 (N2145, N2258);
	BUFX2 g_N2259 (N1000, N2259);
	INVX1 g_N2260 (N3252, N2260);
	INVX1 g_N2261 (N724, N2261);
	BUFX2 g_N2262 (N2588, N2262);
	AND2X1 g_N2263 (N3495, N540, N2263);
	INVX1 g_N2264 (N3635, N2264);
	INVX1 g_N2265 (N3365, N2265);
	INVX1 g_N2266 (N211, N2266);
	INVX1 g_N2267 (N2850, N2267);
	AND2X1 g_N2268 (N3692, N2219, N2268);
	AND2X1 g_N2269 (N200, N90, N2269);
	INVX1 g_N2270 (N161, N2270);
	AND2X1 g_N2271 (N3205, N2837, N2271);
	INVX1 g_N2272 (N503, N2272);
	INVX1 g_N2273 (N2836, N2273);
	INVX1 g_N2274 (N54, N2274);
	INVX1 g_N2275 (N1568, N2275);
	INVX1 g_N2276 (N3355, N2276);
	INVX1 g_N2277 (N132, N2277);
	INVX1 g_N2278 (N1527, N2278);
	AND2X1 g_N2279 (N2067, N3066, N2279);
	INVX1 g_N2280 (N2713, N2280);
	INVX1 g_N2281 (N91, N2281);
	BUFX2 g_N2282 (N2579, N2282);
	INVX1 g_N2283 (N3364, N2283);
	INVX1 g_N2284 (N2216, N2284);
	BUFX2 g_N2285 (N3569, N2285);
	BUFX2 g_N2286 (N2753, N2286);
	BUFX2 g_N321 (N1955, N321);
	INVX1 g_N2287 (N1427, N2287);
	INVX1 g_N2288 (N12, N2288);
	INVX1 g_N2289 (N2706, N2289);
	INVX1 g_N2290 (N256, N2290);
	INVX1 g_N2291 (N3939, N2291);
	AND2X1 g_N2292 (N3097, N515, N2292);
	BUFX2 g_N2293 (N3817, N2293);
	INVX1 g_N2294 (N2859, N2294);
	BUFX2 g_N2295 (N1891, N2295);
	BUFX2 g_N2296 (N3087, N2296);
	INVX1 g_N2297 (N60, N2297);
	INVX1 g_N2298 (N3285, N2298);
	INVX1 g_N2299 (N638, N2299);
	BUFX2 g_N2300 (N1355, N2300);
	AND2X1 g_N2301 (N1708, N3218, N2301);
	INVX1 g_N2302 (N3647, N2302);
	INVX1 g_N2303 (N2097, N2303);
	INVX1 g_N2304 (N124, N2304);
	BUFX2 g_N2305 (N1498, N2305);
	BUFX2 g_N2306 (N3624, N2306);
	BUFX2 g_N2307 (N3744, N2307);
	AND2X1 g_N2308 (N70, N236, N2308);
	BUFX2 g_N2309 (N2401, N2309);
	BUFX2 g_N2310 (N3286, N2310);
	INVX1 g_N2311 (N116, N2311);
	INVX1 g_N2312 (N3764, N2312);
	INVX1 g_N2313 (N1441, N2313);
	BUFX2 g_N2314 (N940, N2314);
	BUFX2 g_N2315 (N3383, N2315);
	BUFX2 g_N2316 (N2918, N2316);
	INVX1 g_N2317 (N1906, N2317);
	BUFX2 g_N2318 (N1594, N2318);
	INVX1 g_N2319 (N53, N2319);
	AND2X1 g_N2320 (N3540, N2111, N2320);
	AND2X1 g_N2321 (N3513, N3173, N2321);
	BUFX2 g_N322 (N458, N322);
	BUFX2 g_N2322 (N3494, N2322);
	AND2X1 g_N2323 (N2463, N3302, N2323);
	AND2X1 g_N2324 (N182, N249, N2324);
	BUFX2 g_N2325 (N3901, N2325);
	AND2X1 g_N2326 (N91, N57, N2326);
	BUFX2 g_N2327 (N3282, N2327);
	INVX1 g_N2328 (N646, N2328);
	BUFX2 g_N2329 (N1961, N2329);
	INVX1 g_N2330 (N487, N2330);
	BUFX2 g_N2331 (N3193, N2331);
	INVX1 g_N2332 (N459, N2332);
	AND2X1 g_N2333 (N2468, N2795, N2333);
	INVX1 g_N2334 (N2932, N2334);
	INVX1 g_N2335 (N231, N2335);
	INVX1 g_N2336 (N3713, N2336);
	BUFX2 g_N2337 (N858, N2337);
	INVX1 g_N2338 (N2719, N2338);
	INVX1 g_N2339 (N140, N2339);
	AND2X1 g_N2340 (N2814, N1546, N2340);
	AND2X1 g_N2341 (N453, N1904, N2341);
	AND2X1 g_N2342 (N2713, N413, N2342);
	AND2X1 g_N2343 (N186, N154, N2343);
	AND2X1 g_N2344 (N2416, N2529, N2344);
	BUFX2 g_N2345 (N3061, N2345);
	AND2X1 g_N2346 (N30, N121, N2346);
	INVX1 g_N2347 (N1013, N2347);
	INVX1 g_N2348 (N3488, N2348);
	BUFX2 g_N2349 (N1438, N2349);
	BUFX2 g_N2350 (N2490, N2350);
	AND2X1 g_N2351 (N3, N226, N2351);
	INVX1 g_N2352 (N902, N2352);
	INVX1 g_N2353 (N246, N2353);
	BUFX2 g_N2354 (N772, N2354);
	INVX1 g_N2355 (N3011, N2355);
	BUFX2 g_N2356 (N2511, N2356);
	INVX1 g_N2357 (N3836, N2357);
	INVX1 g_N2358 (N3393, N2358);
	AND2X1 g_N2359 (N1596, N3369, N2359);
	AND2X1 g_N2360 (N1062, N602, N2360);
	AND2X1 g_N2361 (N203, N63, N2361);
	AND2X1 g_N2362 (N3328, N3425, N2362);
	AND2X1 g_N2363 (N1760, N437, N2363);
	INVX1 g_N2364 (N42, N2364);
	AND2X1 g_N2365 (N3158, N1687, N2365);
	AND2X1 g_N2366 (N3239, N1674, N2366);
	AND2X1 g_N2367 (N153, N99, N2367);
	BUFX2 g_N2368 (N1412, N2368);
	BUFX2 g_N2369 (N3228, N2369);
	AND2X1 g_N2370 (N3204, N1856, N2370);
	BUFX2 g_N2371 (N775, N2371);
	AND2X1 g_N2372 (N1074, N3546, N2372);
	INVX1 g_N2373 (N2924, N2373);
	BUFX2 g_N2374 (N2366, N2374);
	BUFX2 g_N323 (N758, N323);
	INVX1 g_N2375 (N2838, N2375);
	INVX1 g_N2376 (N2494, N2376);
	BUFX2 g_N2377 (N990, N2377);
	BUFX2 g_N2378 (N3572, N2378);
	AND2X1 g_N2379 (N45, N116, N2379);
	BUFX2 g_N2380 (N2916, N2380);
	BUFX2 g_N2381 (N2227, N2381);
	BUFX2 g_N324 (N2153, N324);
	AND2X1 g_N2382 (N2287, N3389, N2382);
	INVX1 g_N2383 (N3272, N2383);
	BUFX2 g_N2384 (N2202, N2384);
	BUFX2 g_N2385 (N2446, N2385);
	INVX1 g_N2386 (N2465, N2386);
	BUFX2 g_N2387 (N3835, N2387);
	BUFX2 g_N2388 (N2006, N2388);
	AND2X1 g_N2389 (N1976, N3876, N2389);
	AND2X1 g_N2390 (N1457, N983, N2390);
	BUFX2 g_N2391 (N2849, N2391);
	INVX1 g_N2392 (N2186, N2392);
	BUFX2 g_N2393 (N3276, N2393);
	BUFX2 g_N2394 (N2652, N2394);
	INVX1 g_N2395 (N1409, N2395);
	INVX1 g_N2396 (N33, N2396);
	INVX1 g_N2397 (N2475, N2397);
	INVX1 g_N2398 (N2859, N2398);
	INVX1 g_N2399 (N1699, N2399);
	BUFX2 g_N2400 (N3568, N2400);
	AND2X1 g_N2401 (N1274, N3109, N2401);
	INVX1 g_N2402 (N534, N2402);
	INVX1 g_N2403 (N1428, N2403);
	BUFX2 g_N2404 (N1239, N2404);
	INVX1 g_N2405 (N201, N2405);
	BUFX2 g_N2406 (N456, N2406);
	INVX1 g_N2407 (N1024, N2407);
	BUFX2 g_N2408 (N1299, N2408);
	INVX1 g_N2409 (N3645, N2409);
	BUFX2 g_N2410 (N401, N2410);
	BUFX2 g_N2411 (N3390, N2411);
	AND2X1 g_N2412 (N656, N1031, N2412);
	BUFX2 g_N2413 (N709, N2413);
	INVX1 g_N2414 (N3931, N2414);
	INVX1 g_N2415 (N1858, N2415);
	BUFX2 g_N2416 (N441, N2416);
	AND2X1 g_N2417 (N3283, N2842, N2417);
	BUFX2 g_N2418 (N1848, N2418);
	INVX1 g_N2419 (N157, N2419);
	BUFX2 g_N2420 (N2874, N2420);
	AND2X1 g_N2421 (N46, N173, N2421);
	INVX1 g_N2422 (N433, N2422);
	AND2X1 g_N2423 (N4, N94, N2423);
	INVX1 g_N2424 (N2737, N2424);
	INVX1 g_N2425 (N2337, N2425);
	INVX1 g_N2426 (N2316, N2426);
	BUFX2 g_N2427 (N2486, N2427);
	INVX1 g_N2428 (N582, N2428);
	BUFX2 g_N2429 (N3769, N2429);
	BUFX2 g_N2430 (N1661, N2430);
	INVX1 g_N2431 (N3303, N2431);
	BUFX2 g_N2432 (N402, N2432);
	BUFX2 g_N2433 (N3435, N2433);
	BUFX2 g_N2434 (N3755, N2434);
	BUFX2 g_N2435 (N3043, N2435);
	INVX1 g_N2436 (N56, N2436);
	BUFX2 g_N325 (N919, N325);
	AND2X1 g_N2437 (N3496, N1413, N2437);
	INVX1 g_N2438 (N2142, N2438);
	INVX1 g_N2439 (N104, N2439);
	INVX1 g_N2440 (N1778, N2440);
	BUFX2 g_N2441 (N1929, N2441);
	AND2X1 g_N2442 (N1157, N1855, N2442);
	INVX1 g_N2443 (N3545, N2443);
	INVX1 g_N2444 (N3886, N2444);
	INVX1 g_N2445 (N2851, N2445);
	AND2X1 g_N2446 (N581, N3032, N2446);
	BUFX2 g_N2447 (N3140, N2447);
	AND2X1 g_N2448 (N386, N2507, N2448);
	AND2X1 g_N2449 (N1484, N2951, N2449);
	AND2X1 g_N2450 (N2698, N3075, N2450);
	AND2X1 g_N2451 (N757, N542, N2451);
	AND2X1 g_N2452 (N3260, N1987, N2452);
	AND2X1 g_N2453 (N799, N1278, N2453);
	BUFX2 g_N326 (N3816, N326);
	INVX1 g_N2454 (N810, N2454);
	AND2X1 g_N2455 (N1263, N3457, N2455);
	BUFX2 g_N2456 (N756, N2456);
	AND2X1 g_N2457 (N1620, N961, N2457);
	INVX1 g_N2458 (N751, N2458);
	AND2X1 g_N2459 (N3046, N2116, N2459);
	AND2X1 g_N2460 (N2626, N1694, N2460);
	INVX1 g_N2461 (N954, N2461);
	INVX1 g_N2462 (N2946, N2462);
	INVX1 g_N2463 (N3195, N2463);
	INVX1 g_N2464 (N501, N2464);
	BUFX2 g_N327 (N1218, N327);
	BUFX2 g_N2465 (N1247, N2465);
	AND2X1 g_N2466 (N2399, N2447, N2466);
	AND2X1 g_N2467 (N2178, N2631, N2467);
	INVX1 g_N2468 (N902, N2468);
	INVX1 g_N2469 (N2257, N2469);
	INVX1 g_N2470 (N1322, N2470);
	INVX1 g_N2471 (N2140, N2471);
	AND2X1 g_N2472 (N1600, N536, N2472);
	BUFX2 g_N2473 (N3007, N2473);
	INVX1 g_N2474 (N2688, N2474);
	BUFX2 g_N2475 (N973, N2475);
	AND2X1 g_N2476 (N1420, N2200, N2476);
	INVX1 g_N2477 (N1030, N2477);
	AND2X1 g_N2478 (N722, N2590, N2478);
	INVX1 g_N2479 (N28, N2479);
	AND2X1 g_N2480 (N3880, N2670, N2480);
	BUFX2 g_N2481 (N1124, N2481);
	AND2X1 g_N2482 (N3313, N2059, N2482);
	INVX1 g_N2483 (N2021, N2483);
	INVX1 g_N2484 (N227, N2484);
	INVX1 g_N2485 (N3434, N2485);
	AND2X1 g_N2486 (N3827, N1677, N2486);
	BUFX2 g_N2487 (N1701, N2487);
	AND2X1 g_N2488 (N3370, N2376, N2488);
	BUFX2 g_N2489 (N3675, N2489);
	AND2X1 g_N2490 (N3474, N981, N2490);
	BUFX2 g_N2491 (N2151, N2491);
	BUFX2 g_N2492 (N2868, N2492);
	BUFX2 g_N2493 (N3671, N2493);
	BUFX2 g_N2494 (N1969, N2494);
	AND2X1 g_N2495 (N41, N169, N2495);
	AND2X1 g_N2496 (N644, N2407, N2496);
	INVX1 g_N2497 (N3355, N2497);
	INVX1 g_N2498 (N3283, N2498);
	AND2X1 g_N2499 (N3210, N2803, N2499);
	BUFX2 g_N2500 (N1560, N2500);
	BUFX2 g_N2501 (N903, N2501);
	AND2X1 g_N2502 (N2177, N1128, N2502);
	BUFX2 g_N2503 (N608, N2503);
	AND2X1 g_N2504 (N2977, N850, N2504);
	INVX1 g_N2505 (N931, N2505);
	BUFX2 g_N2506 (N959, N2506);
	INVX1 g_N2507 (N149, N2507);
	BUFX2 g_N2508 (N1739, N2508);
	BUFX2 g_N2509 (N2892, N2509);
	BUFX2 g_N2510 (N1570, N2510);
	AND2X1 g_N2511 (N3895, N1422, N2511);
	INVX1 g_N2512 (N77, N2512);
	AND2X1 g_N2513 (N3072, N3317, N2513);
	BUFX2 g_N2514 (N777, N2514);
	INVX1 g_N2515 (N2248, N2515);
	AND2X1 g_N2516 (N1726, N2936, N2516);
	INVX1 g_N2517 (N2508, N2517);
	BUFX2 g_N2518 (N680, N2518);
	BUFX2 g_N2519 (N1300, N2519);
	BUFX2 g_N2520 (N3216, N2520);
	AND2X1 g_N2521 (N3900, N2925, N2521);
	INVX1 g_N2522 (N2854, N2522);
	INVX1 g_N2523 (N179, N2523);
	INVX1 g_N2524 (N2706, N2524);
	INVX1 g_N2525 (N1662, N2525);
	INVX1 g_N2526 (N3433, N2526);
	INVX1 g_N2527 (N1084, N2527);
	BUFX2 g_N2528 (N3809, N2528);
	INVX1 g_N2529 (N437, N2529);
	AND2X1 g_N2530 (N1363, N598, N2530);
	BUFX2 g_N2531 (N493, N2531);
	AND2X1 g_N2532 (N972, N1935, N2532);
	INVX1 g_N2533 (N8, N2533);
	INVX1 g_N2534 (N3791, N2534);
	INVX1 g_N2535 (N1402, N2535);
	INVX1 g_N2536 (N79, N2536);
	AND2X1 g_N2537 (N3924, N1553, N2537);
	AND2X1 g_N2538 (N3019, N532, N2538);
	AND2X1 g_N2539 (N498, N3638, N2539);
	BUFX2 g_N2540 (N1669, N2540);
	INVX1 g_N2541 (N1302, N2541);
	BUFX2 g_N2542 (N406, N2542);
	INVX1 g_N2543 (N2187, N2543);
	INVX1 g_N2544 (N847, N2544);
	INVX1 g_N2545 (N2067, N2545);
	AND2X1 g_N2546 (N1314, N828, N2546);
	BUFX2 g_N2547 (N2641, N2547);
	AND2X1 g_N2548 (N3922, N504, N2548);
	AND2X1 g_N2549 (N1605, N2405, N2549);
	BUFX2 g_N2550 (N1352, N2550);
	INVX1 g_N2551 (N2950, N2551);
	INVX1 g_N2552 (N1968, N2552);
	INVX1 g_N2553 (N3242, N2553);
	INVX1 g_N2554 (N1813, N2554);
	AND2X1 g_N2555 (N3113, N3735, N2555);
	INVX1 g_N2556 (N216, N2556);
	AND2X1 g_N2557 (N3294, N1113, N2557);
	INVX1 g_N2558 (N1785, N2558);
	INVX1 g_N2559 (N1748, N2559);
	BUFX2 g_N2560 (N640, N2560);
	BUFX2 g_N2561 (N3366, N2561);
	INVX1 g_N2562 (N677, N2562);
	BUFX2 g_N2563 (N2063, N2563);
	AND2X1 g_N2564 (N2561, N2206, N2564);
	BUFX2 g_N2565 (N1136, N2565);
	AND2X1 g_N2566 (N3509, N1718, N2566);
	INVX1 g_N2567 (N126, N2567);
	BUFX2 g_N2568 (N1860, N2568);
	INVX1 g_N2569 (N1263, N2569);
	BUFX2 g_N2570 (N1939, N2570);
	INVX1 g_N2571 (N152, N2571);
	INVX1 g_N2572 (N6, N2572);
	INVX1 g_N2573 (N3308, N2573);
	INVX1 g_N2574 (N815, N2574);
	AND2X1 g_N2575 (N1384, N1251, N2575);
	BUFX2 g_N2576 (N2450, N2576);
	INVX1 g_N2577 (N1830, N2577);
	AND2X1 g_N2578 (N2358, N3761, N2578);
	AND2X1 g_N2579 (N1913, N2921, N2579);
	AND2X1 g_N2580 (N3887, N3730, N2580);
	BUFX2 g_N2581 (N1626, N2581);
	INVX1 g_N2582 (N3751, N2582);
	INVX1 g_N2583 (N3877, N2583);
	INVX1 g_N2584 (N191, N2584);
	INVX1 g_N2585 (N2138, N2585);
	INVX1 g_N2586 (N2685, N2586);
	INVX1 g_N2587 (N186, N2587);
	AND2X1 g_N2588 (N3068, N1087, N2588);
	AND2X1 g_N2589 (N569, N2643, N2589);
	INVX1 g_N2590 (N1228, N2590);
	AND2X1 g_N2591 (N135, N204, N2591);
	AND2X1 g_N2592 (N1977, N3584, N2592);
	AND2X1 g_N2593 (N535, N3831, N2593);
	INVX1 g_N2594 (N3196, N2594);
	INVX1 g_N2595 (N114, N2595);
	INVX1 g_N2596 (N1194, N2596);
	INVX1 g_N2597 (N2869, N2597);
	BUFX2 g_N328 (N3270, N328);
	AND2X1 g_N2598 (N2220, N2105, N2598);
	BUFX2 g_N2599 (N2549, N2599);
	AND2X1 g_N2600 (N3857, N3740, N2600);
	AND2X1 g_N2601 (N3362, N3038, N2601);
	AND2X1 g_N2602 (N3273, N793, N2602);
	INVX1 g_N2603 (N893, N2603);
	AND2X1 g_N2604 (N2935, N2277, N2604);
	BUFX2 g_N2605 (N695, N2605);
	BUFX2 g_N2606 (N2238, N2606);
	AND2X1 g_N2607 (N3933, N1734, N2607);
	AND2X1 g_N2608 (N3677, N762, N2608);
	BUFX2 g_N2609 (N1348, N2609);
	AND2X1 g_N2610 (N2004, N3056, N2610);
	INVX1 g_N2611 (N3052, N2611);
	INVX1 g_N2612 (N2296, N2612);
	INVX1 g_N2613 (N3491, N2613);
	BUFX2 g_N2614 (N1453, N2614);
	INVX1 g_N2615 (N508, N2615);
	INVX1 g_N2616 (N546, N2616);
	AND2X1 g_N2617 (N2122, N3716, N2617);
	INVX1 g_N2618 (N138, N2618);
	INVX1 g_N2619 (N1684, N2619);
	AND2X1 g_N2620 (N2840, N1959, N2620);
	INVX1 g_N2621 (N184, N2621);
	BUFX2 g_N329 (N1417, N329);
	INVX1 g_N2622 (N1611, N2622);
	BUFX2 g_N2623 (N1184, N2623);
	AND2X1 g_N2624 (N701, N2438, N2624);
	INVX1 g_N2625 (N3339, N2625);
	INVX1 g_N2626 (N178, N2626);
	BUFX2 g_N2627 (N1353, N2627);
	INVX1 g_N2628 (N1, N2628);
	AND2X1 g_N2629 (N3511, N3485, N2629);
	INVX1 g_N2630 (N1868, N2630);
	INVX1 g_N2631 (N1033, N2631);
	AND2X1 g_N2632 (N3632, N1459, N2632);
	INVX1 g_N2633 (N1761, N2633);
	INVX1 g_N2634 (N36, N2634);
	INVX1 g_N2635 (N1235, N2635);
	BUFX2 g_N2636 (N2132, N2636);
	INVX1 g_N2637 (N1913, N2637);
	INVX1 g_N2638 (N3215, N2638);
	BUFX2 g_N2639 (N1604, N2639);
	BUFX2 g_N2640 (N2488, N2640);
	AND2X1 g_N2641 (N3732, N886, N2641);
	BUFX2 g_N2642 (N2229, N2642);
	INVX1 g_N2643 (N2995, N2643);
	BUFX2 g_N2644 (N1951, N2644);
	BUFX2 g_N2645 (N3213, N2645);
	BUFX2 g_N2646 (N3806, N2646);
	BUFX2 g_N2647 (N3264, N2647);
	INVX1 g_N2648 (N1070, N2648);
	AND2X1 g_N2649 (N1451, N1881, N2649);
	BUFX2 g_N2650 (N1650, N2650);
	BUFX2 g_N330 (N818, N330);
	BUFX2 g_N2651 (N3380, N2651);
	AND2X1 g_N2652 (N1489, N1141, N2652);
	BUFX2 g_N2653 (N2039, N2653);
	INVX1 g_N2654 (N2481, N2654);
	AND2X1 g_N2655 (N1103, N1267, N2655);
	BUFX2 g_N2656 (N3665, N2656);
	OR2X1 g_N2657 (N3745, N3119, N2657);
	AND2X1 g_N2658 (N1397, N2523, N2658);
	INVX1 g_N2659 (N2506, N2659);
	BUFX2 g_N2660 (N1117, N2660);
	BUFX2 g_N2661 (N2961, N2661);
	INVX1 g_N2662 (N2100, N2662);
	BUFX2 g_N2663 (N3608, N2663);
	INVX1 g_N2664 (N3302, N2664);
	AND2X1 g_N2665 (N2184, N3181, N2665);
	BUFX2 g_N2666 (N1419, N2666);
	AND2X1 g_N2667 (N1096, N2474, N2667);
	INVX1 g_N2668 (N1168, N2668);
	AND2X1 g_N2669 (N1382, N2087, N2669);
	INVX1 g_N2670 (N73, N2670);
	BUFX2 g_N2671 (N1305, N2671);
	INVX1 g_N2672 (N2209, N2672);
	INVX1 g_N2673 (N1224, N2673);
	INVX1 g_N2674 (N2045, N2674);
	BUFX2 g_N2675 (N3077, N2675);
	INVX1 g_N2676 (N192, N2676);
	INVX1 g_N2677 (N2203, N2677);
	INVX1 g_N2678 (N1607, N2678);
	INVX1 g_N2679 (N2518, N2679);
	AND2X1 g_N2680 (N2891, N2165, N2680);
	INVX1 g_N2681 (N171, N2681);
	AND2X1 g_N2682 (N1454, N1515, N2682);
	AND2X1 g_N2683 (N3152, N837, N2683);
	BUFX2 g_N2684 (N844, N2684);
	BUFX2 g_N2685 (N1308, N2685);
	INVX1 g_N2686 (N776, N2686);
	INVX1 g_N2687 (N100, N2687);
	BUFX2 g_N2688 (N1767, N2688);
	BUFX2 g_N2689 (N398, N2689);
	INVX1 g_N2690 (N2413, N2690);
	INVX1 g_N2691 (N2212, N2691);
	INVX1 g_N2692 (N196, N2692);
	AND2X1 g_N2693 (N120, N89, N2693);
	AND2X1 g_N2694 (N980, N677, N2694);
	INVX1 g_N2695 (N1633, N2695);
	INVX1 g_N2696 (N1954, N2696);
	INVX1 g_N2697 (N2135, N2697);
	INVX1 g_N2698 (N198, N2698);
	BUFX2 g_N2699 (N1823, N2699);
	BUFX2 g_N2700 (N651, N2700);
	BUFX2 g_N2701 (N2459, N2701);
	BUFX2 g_N2702 (N704, N2702);
	AND2X1 g_N2703 (N38, N221, N2703);
	INVX1 g_N2704 (N2660, N2704);
	AND2X1 g_N2705 (N2270, N1789, N2705);
	BUFX2 g_N2706 (N2472, N2706);
	BUFX2 g_N2707 (N3137, N2707);
	INVX1 g_N2708 (N463, N2708);
	AND2X1 g_N2709 (N1916, N1667, N2709);
	AND2X1 g_N2710 (N3284, N488, N2710);
	INVX1 g_N2711 (N3436, N2711);
	AND2X1 g_N2712 (N3566, N3337, N2712);
	BUFX2 g_N2713 (N405, N2713);
	BUFX2 g_N2714 (N1121, N2714);
	INVX1 g_N2715 (N3449, N2715);
	INVX1 g_N2716 (N958, N2716);
	AND2X1 g_N2717 (N241, N37, N2717);
	AND2X1 g_N2718 (N3926, N2414, N2718);
	BUFX2 g_N2719 (N2320, N2719);
	INVX1 g_N2720 (N2209, N2720);
	AND2X1 g_N2721 (N390, N3797, N2721);
	AND2X1 g_N2722 (N3938, N3231, N2722);
	INVX1 g_N2723 (N1517, N2723);
	INVX1 g_N2724 (N1465, N2724);
	INVX1 g_N2725 (N1528, N2725);
	INVX1 g_N2726 (N2154, N2726);
	AND2X1 g_N2727 (N553, N3646, N2727);
	AND2X1 g_N2728 (N3436, N1177, N2728);
	INVX1 g_N2729 (N2198, N2729);
	BUFX2 g_N2730 (N2102, N2730);
	AND2X1 g_N2731 (N513, N3639, N2731);
	AND2X1 g_N2732 (N614, N1794, N2732);
	BUFX2 g_N2733 (N673, N2733);
	AND2X1 g_N2734 (N2280, N3447, N2734);
	INVX1 g_N2735 (N2816, N2735);
	INVX1 g_N2736 (N2286, N2736);
	BUFX2 g_N2737 (N2054, N2737);
	INVX1 g_N2738 (N2305, N2738);
	INVX1 g_N2739 (N3821, N2739);
	BUFX2 g_N2740 (N1245, N2740);
	INVX1 g_N2741 (N1699, N2741);
	INVX1 g_N2742 (N2685, N2742);
	BUFX2 g_N2743 (N3130, N2743);
	BUFX2 g_N2744 (N759, N2744);
	AND2X1 g_N2745 (N3147, N716, N2745);
	INVX1 g_N2746 (N481, N2746);
	BUFX2 g_N2747 (N2997, N2747);
	BUFX2 g_N2748 (N1236, N2748);
	BUFX2 g_N2749 (N1938, N2749);
	AND2X1 g_N2750 (N219, N108, N2750);
	INVX1 g_N2751 (N61, N2751);
	BUFX2 g_N2752 (N485, N2752);
	AND2X1 g_N2753 (N928, N3131, N2753);
	BUFX2 g_N2754 (N2096, N2754);
	AND2X1 g_N2755 (N223, N193, N2755);
	BUFX2 g_N2756 (N489, N2756);
	INVX1 g_N2757 (N760, N2757);
	BUFX2 g_N2758 (N1371, N2758);
	INVX1 g_N2759 (N649, N2759);
	AND2X1 g_N2760 (N1803, N1706, N2760);
	INVX1 g_N2761 (N3198, N2761);
	AND2X1 g_N2762 (N1984, N2160, N2762);
	AND2X1 g_N2763 (N1473, N1035, N2763);
	INVX1 g_N2764 (N1744, N2764);
	INVX1 g_N2765 (N172, N2765);
	INVX1 g_N2766 (N930, N2766);
	BUFX2 g_N2767 (N1321, N2767);
	AND2X1 g_N2768 (N2986, N3157, N2768);
	INVX1 g_N2769 (N2831, N2769);
	INVX1 g_N2770 (N2109, N2770);
	BUFX2 g_N2771 (N1106, N2771);
	INVX1 g_N2772 (N3407, N2772);
	INVX1 g_N2773 (N222, N2773);
	INVX1 g_N2774 (N253, N2774);
	INVX1 g_N2775 (N2864, N2775);
	INVX1 g_N2776 (N1645, N2776);
	INVX1 g_N2777 (N3298, N2777);
	INVX1 g_N2778 (N1480, N2778);
	INVX1 g_N2779 (N2914, N2779);
	AND2X1 g_N2780 (N115, N155, N2780);
	BUFX2 g_N2781 (N477, N2781);
	AND2X1 g_N2782 (N1212, N969, N2782);
	INVX1 g_N2783 (N235, N2783);
	BUFX2 g_N2784 (N3145, N2784);
	BUFX2 g_N2785 (N3412, N2785);
	INVX1 g_N2786 (N2349, N2786);
	AND2X1 g_N2787 (N2112, N2800, N2787);
	INVX1 g_N2788 (N2945, N2788);
	AND2X1 g_N2789 (N1817, N2587, N2789);
	AND2X1 g_N2790 (N942, N1206, N2790);
	INVX1 g_N2791 (N3543, N2791);
	AND2X1 g_N2792 (N1001, N1100, N2792);
	INVX1 g_N2793 (N141, N2793);
	INVX1 g_N2794 (N48, N2794);
	INVX1 g_N2795 (N2550, N2795);
	AND2X1 g_N2796 (N708, N1962, N2796);
	AND2X1 g_N2797 (N2431, N1567, N2797);
	BUFX2 g_N2798 (N1038, N2798);
	INVX1 g_N2799 (N846, N2799);
	INVX1 g_N2800 (N2354, N2800);
	INVX1 g_N2801 (N1084, N2801);
	INVX1 g_N2802 (N2078, N2802);
	INVX1 g_N2803 (N2300, N2803);
	INVX1 g_N2804 (N479, N2804);
	INVX1 g_N2805 (N2236, N2805);
	BUFX2 g_N2806 (N3890, N2806);
	BUFX2 g_N2807 (N932, N2807);
	INVX1 g_N2808 (N3447, N2808);
	BUFX2 g_N2809 (N3445, N2809);
	BUFX2 g_N2810 (N1110, N2810);
	BUFX2 g_N2811 (N1814, N2811);
	INVX1 g_N2812 (N1221, N2812);
	BUFX2 g_N2813 (N2601, N2813);
	INVX1 g_N2814 (N2356, N2814);
	AND2X1 g_N2815 (N111, N244, N2815);
	BUFX2 g_N2816 (N3514, N2816);
	INVX1 g_N2817 (N203, N2817);
	AND2X1 g_N2818 (N2256, N1712, N2818);
	INVX1 g_N2819 (N3235, N2819);
	AND2X1 g_N2820 (N1200, N1627, N2820);
	AND2X1 g_N2821 (N1610, N1185, N2821);
	AND2X1 g_N2822 (N571, N3724, N2822);
	AND2X1 g_N2823 (N2966, N874, N2823);
	AND2X1 g_N2824 (N1223, N3609, N2824);
	AND2X1 g_N2825 (N1736, N2477, N2825);
	AND2X1 g_N2826 (N2970, N1614, N2826);
	BUFX2 g_N2827 (N1577, N2827);
	AND2X1 g_N2828 (N3497, N1302, N2828);
	INVX1 g_N2829 (N3194, N2829);
	INVX1 g_N2830 (N1055, N2830);
	BUFX2 g_N2831 (N3004, N2831);
	INVX1 g_N2832 (N30, N2832);
	INVX1 g_N2833 (N862, N2833);
	BUFX2 g_N2834 (N854, N2834);
	INVX1 g_N2835 (N2152, N2835);
	BUFX2 g_N2836 (N3760, N2836);
	INVX1 g_N2837 (N2394, N2837);
	BUFX2 g_N2838 (N3768, N2838);
	INVX1 g_N2839 (N2249, N2839);
	INVX1 g_N2840 (N23, N2840);
	AND2X1 g_N2841 (N3025, N1625, N2841);
	INVX1 g_N2842 (N987, N2842);
	AND2X1 g_N2843 (N2373, N1583, N2843);
	INVX1 g_N2844 (N2899, N2844);
	BUFX2 g_N2845 (N2323, N2845);
	INVX1 g_N2846 (N690, N2846);
	INVX1 g_N2847 (N1046, N2847);
	BUFX2 g_N2848 (N925, N2848);
	AND2X1 g_N2849 (N2786, N2672, N2849);
	BUFX2 g_N2850 (N1208, N2850);
	BUFX2 g_N2851 (N3757, N2851);
	INVX1 g_N2852 (N425, N2852);
	AND2X1 g_N2853 (N2863, N1875, N2853);
	BUFX2 g_N2854 (N624, N2854);
	BUFX2 g_N2855 (N1166, N2855);
	INVX1 g_N2856 (N1763, N2856);
	INVX1 g_N2857 (N870, N2857);
	BUFX2 g_N2858 (N3084, N2858);
	BUFX2 g_N2859 (N1808, N2859);
	BUFX2 g_N2860 (N1209, N2860);
	BUFX2 g_N2861 (N1080, N2861);
	INVX1 g_N2862 (N699, N2862);
	INVX1 g_N2863 (N391, N2863);
	BUFX2 g_N2864 (N3168, N2864);
	INVX1 g_N2865 (N3699, N2865);
	AND2X1 g_N2866 (N993, N3582, N2866);
	AND2X1 g_N2867 (N3138, N830, N2867);
	AND2X1 g_N2868 (N47, N180, N2868);
	BUFX2 g_N2869 (N3414, N2869);
	BUFX2 g_N2870 (N3050, N2870);
	AND2X1 g_N2871 (N1181, N1279, N2871);
	INVX1 g_N2872 (N237, N2872);
	INVX1 g_N2873 (N2080, N2873);
	AND2X1 g_N2874 (N2716, N3770, N2874);
	BUFX2 g_N2875 (N1172, N2875);
	AND2X1 g_N2876 (N597, N1721, N2876);
	BUFX2 g_N2877 (N3679, N2877);
	AND2X1 g_N2878 (N3935, N804, N2878);
	INVX1 g_N2879 (N144, N2879);
	AND2X1 g_N2880 (N2353, N2765, N2880);
	AND2X1 g_N2881 (N2621, N1963, N2881);
	AND2X1 g_N2882 (N2338, N502, N2882);
	BUFX2 g_N331 (N3541, N331);
	AND2X1 g_N2883 (N688, N3030, N2883);
	INVX1 g_N2884 (N3437, N2884);
	AND2X1 g_N2885 (N2933, N2015, N2885);
	INVX1 g_N2886 (N2642, N2886);
	INVX1 g_N2887 (N3629, N2887);
	INVX1 g_N2888 (N875, N2888);
	BUFX2 g_N2889 (N3462, N2889);
	INVX1 g_N2890 (N2831, N2890);
	INVX1 g_N2891 (N1746, N2891);
	AND2X1 g_N2892 (N2335, N451, N2892);
	INVX1 g_N2893 (N1343, N2893);
	BUFX2 g_N2894 (N1368, N2894);
	BUFX2 g_N2895 (N3879, N2895);
	AND2X1 g_N2896 (N1163, N2662, N2896);
	BUFX2 g_N332 (N464, N332);
	AND2X1 g_N2897 (N3941, N2615, N2897);
	BUFX2 g_N333 (N1958, N333);
	INVX1 g_N2898 (N778, N2898);
	BUFX2 g_N2899 (N3525, N2899);
	INVX1 g_N2900 (N1967, N2900);
	AND2X1 g_N2901 (N2226, N1649, N2901);
	BUFX2 g_N2902 (N1383, N2902);
	BUFX2 g_N2903 (N842, N2903);
	INVX1 g_N2904 (N51, N2904);
	BUFX2 g_N334 (N3583, N334);
	AND2X1 g_N2905 (N71, N93, N2905);
	AND2X1 g_N2906 (N1840, N1755, N2906);
	AND2X1 g_N2907 (N3862, N3002, N2907);
	INVX1 g_N2908 (N156, N2908);
	INVX1 g_N2909 (N953, N2909);
	INVX1 g_N2910 (N827, N2910);
	AND2X1 g_N2911 (N881, N924, N2911);
	AND2X1 g_N2912 (N1388, N2355, N2912);
	INVX1 g_N2913 (N496, N2913);
	BUFX2 g_N2914 (N2649, N2914);
	BUFX2 g_N335 (N1174, N335);
	AND2X1 g_N2915 (N243, N124, N2915);
	AND2X1 g_N2916 (N3908, N668, N2916);
	AND2X1 g_N2917 (N3787, N1349, N2917);
	AND2X1 g_N2918 (N1532, N2487, N2918);
	AND2X1 g_N2919 (N814, N719, N2919);
	BUFX2 g_N2920 (N3907, N2920);
	INVX1 g_N2921 (N1310, N2921);
	BUFX2 g_N2922 (N897, N2922);
	INVX1 g_N2923 (N3535, N2923);
	BUFX2 g_N2924 (N2361, N2924);
	INVX1 g_N2925 (N884, N2925);
	BUFX2 g_N2926 (N2843, N2926);
	BUFX2 g_N2927 (N3340, N2927);
	AND2X1 g_N2928 (N2290, N429, N2928);
	INVX1 g_N2929 (N1041, N2929);
	AND2X1 g_N2930 (N131, N170, N2930);
	BUFX2 g_N336 (N3779, N336);
	BUFX2 g_N2931 (N2128, N2931);
	BUFX2 g_N2932 (N1292, N2932);
	BUFX2 g_N337 (N2307, N337);
	BUFX2 g_N2933 (N1776, N2933);
	AND2X1 g_N2934 (N1306, N1408, N2934);
	INVX1 g_N2935 (N62, N2935);
	INVX1 g_N2936 (N1811, N2936);
	AND2X1 g_N2937 (N3789, N3154, N2937);
	INVX1 g_N2938 (N2035, N2938);
	BUFX2 g_N2939 (N2591, N2939);
	BUFX2 g_N2940 (N3429, N2940);
	INVX1 g_N2941 (N2388, N2941);
	INVX1 g_N2942 (N3564, N2942);
	AND2X1 g_N2943 (N139, N2, N2943);
	INVX1 g_N2944 (N3478, N2944);
	BUFX2 g_N2945 (N3763, N2945);
	BUFX2 g_N2946 (N785, N2946);
	AND2X1 g_N2947 (N1732, N2107, N2947);
	BUFX2 g_N2948 (N3602, N2948);
	INVX1 g_N2949 (N534, N2949);
	BUFX2 g_N2950 (N3301, N2950);
	BUFX2 g_N2951 (N3310, N2951);
	BUFX2 g_N2952 (N2346, N2952);
	INVX1 g_N2953 (N2933, N2953);
	INVX1 g_N2954 (N649, N2954);
	INVX1 g_N2955 (N3303, N2955);
	INVX1 g_N2956 (N2146, N2956);
	INVX1 g_N2957 (N2207, N2957);
	INVX1 g_N2958 (N1327, N2958);
	AND2X1 g_N2959 (N936, N1376, N2959);
	BUFX2 g_N2960 (N3034, N2960);
	AND2X1 g_N2961 (N183, N100, N2961);
	AND2X1 g_N2962 (N9, N137, N2962);
	AND2X1 g_N2963 (N16, N237, N2963);
	BUFX2 g_N2964 (N3081, N2964);
	INVX1 g_N2965 (N1047, N2965);
	INVX1 g_N2966 (N2964, N2966);
	BUFX2 g_N338 (N444, N338);
	BUFX2 g_N2967 (N2333, N2967);
	INVX1 g_N2968 (N3368, N2968);
	INVX1 g_N2969 (N2215, N2969);
	INVX1 g_N2970 (N74, N2970);
	INVX1 g_N2971 (N914, N2971);
	INVX1 g_N2972 (N3402, N2972);
	INVX1 g_N2973 (N234, N2973);
	BUFX2 g_N2974 (N3618, N2974);
	BUFX2 g_N2975 (N1447, N2975);
	BUFX2 g_N2976 (N1054, N2976);
	INVX1 g_N2977 (N3327, N2977);
	INVX1 g_N2978 (N1328, N2978);
	AND2X1 g_N2979 (N438, N3451, N2979);
	INVX1 g_N2980 (N2903, N2980);
	BUFX2 g_N2981 (N440, N2981);
	AND2X1 g_N2982 (N2289, N1098, N2982);
	INVX1 g_N2983 (N1813, N2983);
	INVX1 g_N2984 (N3594, N2984);
	INVX1 g_N2985 (N3422, N2985);
	INVX1 g_N2986 (N1466, N2986);
	AND2X1 g_N2987 (N1164, N2847, N2987);
	AND2X1 g_N2988 (N2021, N832, N2988);
	INVX1 g_N2989 (N3906, N2989);
	INVX1 g_N2990 (N958, N2990);
	INVX1 g_N2991 (N3419, N2991);
	BUFX2 g_N2992 (N2342, N2992);
	AND2X1 g_N2993 (N166, N143, N2993);
	INVX1 g_N2994 (N1027, N2994);
	BUFX2 g_N2995 (N1012, N2995);
	INVX1 g_N2996 (N1329, N2996);
	AND2X1 g_N2997 (N2180, N3854, N2997);
	AND2X1 g_N2998 (N2368, N2386, N2998);
	INVX1 g_N2999 (N2371, N2999);
	INVX1 g_N3000 (N2137, N3000);
	INVX1 g_N3001 (N188, N3001);
	INVX1 g_N3002 (N1742, N3002);
	BUFX2 g_N3003 (N1666, N3003);
	AND2X1 g_N3004 (N2739, N2696, N3004);
	INVX1 g_N3005 (N773, N3005);
	AND2X1 g_N3006 (N491, N3774, N3006);
	AND2X1 g_N3007 (N422, N1552, N3007);
	INVX1 g_N3008 (N1906, N3008);
	INVX1 g_N3009 (N3591, N3009);
	BUFX2 g_N3010 (N939, N3010);
	BUFX2 g_N339 (N3912, N339);
	BUFX2 g_N3011 (N3921, N3011);
	INVX1 g_N3012 (N47, N3012);
	INVX1 g_N3013 (N2663, N3013);
	INVX1 g_N3014 (N1333, N3014);
	BUFX2 g_N3015 (N833, N3015);
	AND2X1 g_N3016 (N1558, N3942, N3016);
	AND2X1 g_N3017 (N246, N172, N3017);
	BUFX2 g_N3018 (N1145, N3018);
	INVX1 g_N3019 (N199, N3019);
	INVX1 g_N3020 (N3141, N3020);
	AND2X1 g_N3021 (N1565, N3175, N3021);
	INVX1 g_N3022 (N2974, N3022);
	INVX1 g_N3023 (N107, N3023);
	INVX1 g_N3024 (N3906, N3024);
	INVX1 g_N3025 (N11, N3025);
	AND2X1 g_N3026 (N1226, N1341, N3026);
	AND2X1 g_N3027 (N3529, N3365, N3027);
	INVX1 g_N3028 (N2019, N3028);
	INVX1 g_N3029 (N3260, N3029);
	INVX1 g_N3030 (N578, N3030);
	INVX1 g_N3031 (N3656, N3031);
	INVX1 g_N3032 (N1491, N3032);
	BUFX2 g_N3033 (N3533, N3033);
	AND2X1 g_N3034 (N3319, N664, N3034);
	BUFX2 g_N3035 (N1264, N3035);
	BUFX2 g_N3036 (N1887, N3036);
	BUFX2 g_N3037 (N1463, N3037);
	INVX1 g_N3038 (N888, N3038);
	INVX1 g_N3039 (N459, N3039);
	INVX1 g_N3040 (N476, N3040);
	INVX1 g_N3041 (N1575, N3041);
	INVX1 g_N3042 (N3436, N3042);
	AND2X1 g_N3043 (N2328, N591, N3043);
	INVX1 g_N3044 (N57, N3044);
	INVX1 g_N3045 (N589, N3045);
	INVX1 g_N3046 (N824, N3046);
	INVX1 g_N3047 (N796, N3047);
	INVX1 g_N3048 (N3356, N3048);
	AND2X1 g_N3049 (N1869, N1486, N3049);
	AND2X1 g_N3050 (N39, N32, N3050);
	BUFX2 g_N3051 (N1543, N3051);
	BUFX2 g_N3052 (N3683, N3052);
	INVX1 g_N3053 (N3502, N3053);
	BUFX2 g_N3054 (N3704, N3054);
	BUFX2 g_N3055 (N1937, N3055);
	INVX1 g_N3056 (N110, N3056);
	BUFX2 g_N3057 (N1928, N3057);
	BUFX2 g_N340 (N3614, N340);
	BUFX2 g_N3058 (N819, N3058);
	BUFX2 g_N3059 (N744, N3059);
	INVX1 g_N3060 (N1083, N3060);
	AND2X1 g_N3061 (N2788, N3604, N3061);
	INVX1 g_N3062 (N494, N3062);
	BUFX2 g_N3063 (N2911, N3063);
	INVX1 g_N3064 (N1342, N3064);
	AND2X1 g_N3065 (N901, N2677, N3065);
	INVX1 g_N3066 (N1873, N3066);
	AND2X1 g_N3067 (N3316, N2612, N3067);
	INVX1 g_N3068 (N566, N3068);
	BUFX2 g_N3069 (N2912, N3069);
	BUFX2 g_N3070 (N2709, N3070);
	BUFX2 g_N3071 (N2029, N3071);
	INVX1 g_N3072 (N889, N3072);
	AND2X1 g_N3073 (N3810, N3651, N3073);
	INVX1 g_N3074 (N3916, N3074);
	INVX1 g_N3075 (N230, N3075);
	AND2X1 g_N3076 (N2398, N2246, N3076);
	AND2X1 g_N3077 (N2715, N2175, N3077);
	BUFX2 g_N3078 (N650, N3078);
	AND2X1 g_N3079 (N2284, N3295, N3079);
	BUFX2 g_N3080 (N845, N3080);
	AND2X1 g_N3081 (N3673, N394, N3081);
	BUFX2 g_N3082 (N2928, N3082);
	AND2X1 g_N3083 (N3208, N3893, N3083);
	AND2X1 g_N3084 (N17, N175, N3084);
	AND2X1 g_N3085 (N1049, N1588, N3085);
	BUFX2 g_N3086 (N2792, N3086);
	AND2X1 g_N3087 (N555, N3169, N3087);
	BUFX2 g_N3088 (N3162, N3088);
	AND2X1 g_N3089 (N3838, N3118, N3089);
	INVX1 g_N3090 (N3939, N3090);
	AND2X1 g_N3091 (N3731, N2066, N3091);
	INVX1 g_N3092 (N2902, N3092);
	BUFX2 g_N3093 (N866, N3093);
	BUFX2 g_N3094 (N3126, N3094);
	INVX1 g_N3095 (N739, N3095);
	AND2X1 g_N3096 (N3028, N1242, N3096);
	INVX1 g_N3097 (N1470, N3097);
	INVX1 g_N3098 (N1621, N3098);
	INVX1 g_N3099 (N798, N3099);
	INVX1 g_N3100 (N40, N3100);
	AND2X1 g_N3101 (N3824, N3520, N3101);
	BUFX2 g_N341 (N3315, N341);
	INVX1 g_N3102 (N2131, N3102);
	INVX1 g_N3103 (N3253, N3103);
	INVX1 g_N3104 (N966, N3104);
	INVX1 g_N3105 (N1395, N3105);
	AND2X1 g_N3106 (N1290, N3512, N3106);
	INVX1 g_N3107 (N1742, N3107);
	INVX1 g_N3108 (N1440, N3108);
	INVX1 g_N3109 (N3058, N3109);
	BUFX2 g_N3110 (N1186, N3110);
	INVX1 g_N3111 (N1838, N3111);
	INVX1 g_N3112 (N135, N3112);
	INVX1 g_N3113 (N217, N3113);
	INVX1 g_N3114 (N1872, N3114);
	AND2X1 g_N3115 (N3833, N3246, N3115);
	INVX1 g_N3116 (N3807, N3116);
	BUFX2 g_N3117 (N1332, N3117);
	INVX1 g_N3118 (N2349, N3118);
	BUFX2 g_N3119 (N1253, N3119);
	AND2X1 g_N3120 (N3670, N3657, N3120);
	AND2X1 g_N3121 (N110, N220, N3121);
	AND2X1 g_N3122 (N460, N3689, N3122);
	AND2X1 g_N3123 (N2443, N1203, N3123);
	INVX1 g_N3124 (N2212, N3124);
	INVX1 g_N3125 (N1295, N3125);
	AND2X1 g_N3126 (N2938, N3350, N3126);
	AND2X1 g_N3127 (N1120, N1864, N3127);
	INVX1 g_N3128 (N642, N3128);
	BUFX2 g_N342 (N3086, N342);
	BUFX2 g_N3129 (N2379, N3129);
	AND2X1 g_N3130 (N15, N127, N3130);
	INVX1 g_N3131 (N1682, N3131);
	BUFX2 g_N343 (N3010, N343);
	INVX1 g_N3132 (N1450, N3132);
	AND2X1 g_N3133 (N27, N196, N3133);
	INVX1 g_N3134 (N2700, N3134);
	INVX1 g_N3135 (N1435, N3135);
	INVX1 g_N3136 (N239, N3136);
	AND2X1 g_N3137 (N3220, N745, N3137);
	INVX1 g_N3138 (N3938, N3138);
	INVX1 g_N3139 (N3673, N3139);
	AND2X1 g_N3140 (N1456, N3114, N3140);
	BUFX2 g_N3141 (N3049, N3141);
	BUFX2 g_N3142 (N1469, N3142);
	BUFX2 g_N3143 (N2905, N3143);
	INVX1 g_N3144 (N2447, N3144);
	AND2X1 g_N3145 (N2278, N2422, N3145);
	INVX1 g_N3146 (N3524, N3146);
	INVX1 g_N3147 (N3739, N3147);
	INVX1 g_N3148 (N929, N3148);
	BUFX2 g_N3149 (N3709, N3149);
	BUFX2 g_N344 (N3871, N344);
	BUFX2 g_N3150 (N2012, N3150);
	INVX1 g_N3151 (N1006, N3151);
	INVX1 g_N3152 (N3636, N3152);
	BUFX2 g_N345 (N400, N345);
	INVX1 g_N3153 (N2976, N3153);
	INVX1 g_N3154 (N19, N3154);
	AND2X1 g_N3155 (N1638, N1990, N3155);
	BUFX2 g_N3156 (N556, N3156);
	INVX1 g_N3157 (N2186, N3157);
	INVX1 g_N3158 (N2568, N3158);
	AND2X1 g_N3159 (N1953, N3100, N3159);
	INVX1 g_N3160 (N2296, N3160);
	AND2X1 g_N3161 (N82, N21, N3161);
	AND2X1 g_N3162 (N1949, N1585, N3162);
	INVX1 g_N3163 (N1278, N3163);
	INVX1 g_N3164 (N1343, N3164);
	BUFX2 g_N3165 (N3856, N3165);
	INVX1 g_N3166 (N1819, N3166);
	AND2X1 g_N3167 (N548, N2117, N3167);
	BUFX2 g_N346 (N2181, N346);
	AND2X1 g_N3168 (N1435, N2844, N3168);
	INVX1 g_N3169 (N214, N3169);
	AND2X1 g_N3170 (N1483, N1060, N3170);
	INVX1 g_N3171 (N3491, N3171);
	INVX1 g_N3172 (N2020, N3172);
	INVX1 g_N3173 (N173, N3173);
	INVX1 g_N3174 (N3365, N3174);
	INVX1 g_N3175 (N481, N3175);
	INVX1 g_N3176 (N183, N3176);
	BUFX2 g_N347 (N3888, N347);
	INVX1 g_N3177 (N550, N3177);
	AND2X1 g_N3178 (N2262, N1643, N3178);
	INVX1 g_N3179 (N109, N3179);
	AND2X1 g_N3180 (N2242, N2000, N3180);
	INVX1 g_N3181 (N3627, N3181);
	AND2X1 g_N3182 (N1601, N2043, N3182);
	INVX1 g_N3183 (N773, N3183);
	BUFX2 g_N348 (N3377, N348);
	INVX1 g_N3184 (N166, N3184);
	INVX1 g_N3185 (N247, N3185);
	AND2X1 g_N3186 (N672, N2298, N3186);
	AND2X1 g_N3187 (N3686, N2265, N3187);
	AND2X1 g_N3188 (N2215, N1088, N3188);
	AND2X1 g_N3189 (N2770, N1657, N3189);
	BUFX2 g_N3190 (N643, N3190);
	BUFX2 g_N3191 (N1132, N3191);
	BUFX2 g_N3192 (N1439, N3192);
	AND2X1 g_N3193 (N114, N148, N3193);
	BUFX2 g_N3194 (N1934, N3194);
	BUFX2 g_N3195 (N1702, N3195);
	BUFX2 g_N3196 (N2790, N3196);
	AND2X1 g_N3197 (N472, N447, N3197);
	BUFX2 g_N3198 (N1125, N3198);
	AND2X1 g_N3199 (N884, N1564, N3199);
	BUFX2 g_N3200 (N2011, N3200);
	INVX1 g_N3201 (N3540, N3201);
	INVX1 g_N3202 (N2889, N3202);
	AND2X1 g_N3203 (N2950, N593, N3203);
	INVX1 g_N3204 (N2156, N3204);
	BUFX2 g_N3205 (N1072, N3205);
	AND2X1 g_N3206 (N2533, N2244, N3206);
	BUFX2 g_N3207 (N3256, N3207);
	INVX1 g_N3208 (N1010, N3208);
	AND2X1 g_N3209 (N3334, N3615, N3209);
	INVX1 g_N3210 (N408, N3210);
	BUFX2 g_N3211 (N2451, N3211);
	INVX1 g_N3212 (N2606, N3212);
	AND2X1 g_N3213 (N1973, N1499, N3213);
	INVX1 g_N3214 (N1077, N3214);
	BUFX2 g_N349 (N666, N349);
	BUFX2 g_N3215 (N3324, N3215);
	AND2X1 g_N3216 (N2996, N1445, N3216);
	BUFX2 g_N3217 (N2163, N3217);
	INVX1 g_N3218 (N3337, N3218);
	INVX1 g_N3219 (N202, N3219);
	INVX1 g_N3220 (N746, N3220);
	AND2X1 g_N3221 (N199, N145, N3221);
	INVX1 g_N3222 (N439, N3222);
	BUFX2 g_N3223 (N592, N3223);
	AND2X1 g_N3224 (N2055, N1241, N3224);
	BUFX2 g_N350 (N1787, N350);
	BUFX2 g_N3225 (N2694, N3225);
	INVX1 g_N3226 (N3717, N3226);
	BUFX2 g_N351 (N805, N351);
	AND2X1 g_N3227 (N1908, N1968, N3227);
	AND2X1 g_N3228 (N3299, N2394, N3228);
	INVX1 g_N3229 (N1237, N3229);
	AND2X1 g_N3230 (N611, N3080, N3230);
	INVX1 g_N3231 (N1982, N3231);
	INVX1 g_N3232 (N1224, N3232);
	INVX1 g_N3233 (N2570, N3233);
	INVX1 g_N3234 (N976, N3234);
	BUFX2 g_N3235 (N3360, N3235);
	INVX1 g_N3236 (N2875, N3236);
	BUFX2 g_N3237 (N1673, N3237);
	BUFX2 g_N3238 (N1723, N3238);
	INVX1 g_N3239 (N2441, N3239);
	AND2X1 g_N3240 (N648, N1131, N3240);
	INVX1 g_N3241 (N1062, N3241);
	BUFX2 g_N3242 (N3209, N3242);
	AND2X1 g_N3243 (N3283, N1105, N3243);
	AND2X1 g_N3244 (N3132, N2309, N3244);
	AND2X1 g_N3245 (N2525, N642, N3245);
	INVX1 g_N3246 (N3312, N3246);
	AND2X1 g_N3247 (N3196, N560, N3247);
	INVX1 g_N3248 (N764, N3248);
	INVX1 g_N3249 (N1933, N3249);
	INVX1 g_N3250 (N3635, N3250);
	INVX1 g_N3251 (N3420, N3251);
	BUFX2 g_N3252 (N2937, N3252);
	BUFX2 g_N3253 (N1644, N3253);
	BUFX2 g_N3254 (N2245, N3254);
	INVX1 g_N3255 (N3367, N3255);
	BUFX2 g_N352 (N2975, N352);
	AND2X1 g_N3256 (N637, N3306, N3256);
	AND2X1 g_N3257 (N392, N465, N3257);
	BUFX2 g_N3258 (N1115, N3258);
	INVX1 g_N3259 (N2542, N3259);
	BUFX2 g_N3260 (N2390, N3260);
	AND2X1 g_N3261 (N776, N2336, N3261);
	INVX1 g_N3262 (N3143, N3262);
	AND2X1 g_N3263 (N3185, N2266, N3263);
	AND2X1 g_N3264 (N915, N1672, N3264);
	INVX1 g_N3265 (N1082, N3265);
	INVX1 g_N3266 (N2385, N3266);
	INVX1 g_N3267 (N139, N3267);
	BUFX2 g_N3268 (N774, N3268);
	BUFX2 g_N3269 (N1749, N3269);
	BUFX2 g_N3270 (N480, N3270);
	BUFX2 g_N353 (N3841, N353);
	INVX1 g_N3271 (N1549, N3271);
	BUFX2 g_N3272 (N1985, N3272);
	INVX1 g_N3273 (N190, N3273);
	INVX1 g_N3274 (N1448, N3274);
	INVX1 g_N3275 (N3371, N3275);
	AND2X1 g_N3276 (N1432, N1613, N3276);
	BUFX2 g_N3277 (N3159, N3277);
	INVX1 g_N3278 (N3588, N3278);
	BUFX2 g_N3279 (N1381, N3279);
	BUFX2 g_N3280 (N557, N3280);
	INVX1 g_N3281 (N3191, N3281);
	AND2X1 g_N3282 (N3711, N1370, N3282);
	BUFX2 g_N3283 (N2324, N3283);
	INVX1 g_N3284 (N193, N3284);
	BUFX2 g_N3285 (N1563, N3285);
	AND2X1 g_N3286 (N1108, N2766, N3286);
	AND2X1 g_N3287 (N3172, N1244, N3287);
	BUFX2 g_N3288 (N1366, N3288);
	AND2X1 g_N3289 (N2176, N2275, N3289);
	INVX1 g_N3290 (N3927, N3290);
	INVX1 g_N3291 (N2858, N3291);
	BUFX2 g_N3292 (N3904, N3292);
	BUFX2 g_N3293 (N3188, N3293);
	BUFX2 g_N354 (N2771, N354);
	INVX1 g_N3294 (N1983, N3294);
	INVX1 g_N3295 (N1980, N3295);
	INVX1 g_N3296 (N1410, N3296);
	AND2X1 g_N3297 (N2375, N1740, N3297);
	BUFX2 g_N3298 (N1032, N3298);
	INVX1 g_N3299 (N3205, N3299);
	INVX1 g_N3300 (N241, N3300);
	AND2X1 g_N3301 (N3650, N3212, N3301);
	BUFX2 g_N3302 (N3516, N3302);
	BUFX2 g_N3303 (N2555, N3303);
	BUFX2 g_N3304 (N3320, N3304);
	INVX1 g_N3305 (N1772, N3305);
	INVX1 g_N3306 (N601, N3306);
	AND2X1 g_N3307 (N1629, N2364, N3307);
	BUFX2 g_N3308 (N2680, N3308);
	INVX1 g_N3309 (N1691, N3309);
	AND2X1 g_N3310 (N3399, N1173, N3310);
	BUFX2 g_N3311 (N906, N3311);
	BUFX2 g_N3312 (N1795, N3312);
	INVX1 g_N3313 (N628, N3313);
	BUFX2 g_N3314 (N734, N3314);
	BUFX2 g_N3315 (N1019, N3315);
	INVX1 g_N3316 (N3198, N3316);
	INVX1 g_N3317 (N2920, N3317);
	AND2X1 g_N3318 (N3902, N2551, N3318);
	BUFX2 g_N355 (N1429, N355);
	INVX1 g_N3319 (N18, N3319);
	AND2X1 g_N3320 (N2900, N2802, N3320);
	AND2X1 g_N3321 (N2193, N1283, N3321);
	BUFX2 g_N3322 (N1874, N3322);
	INVX1 g_N3323 (N1914, N3323);
	AND2X1 g_N3324 (N2835, N1773, N3324);
	INVX1 g_N3325 (N2240, N3325);
	INVX1 g_N3326 (N2748, N3326);
	BUFX2 g_N3327 (N3820, N3327);
	INVX1 g_N3328 (N1416, N3328);
	INVX1 g_N3329 (N2636, N3329);
	BUFX2 g_N3330 (N736, N3330);
	AND2X1 g_N3331 (N872, N3633, N3331);
	BUFX2 g_N3332 (N544, N3332);
	INVX1 g_N3333 (N2080, N3333);
	INVX1 g_N3334 (N3782, N3334);
	BUFX2 g_N3335 (N1323, N3335);
	BUFX2 g_N3336 (N2598, N3336);
	BUFX2 g_N3337 (N2197, N3337);
	AND2X1 g_N3338 (N654, N2069, N3338);
	BUFX2 g_N356 (N2038, N356);
	BUFX2 g_N3339 (N1029, N3339);
	AND2X1 g_N3340 (N3778, N2313, N3340);
	INVX1 g_N3341 (N3595, N3341);
	AND2X1 g_N3342 (N1482, N3934, N3342);
	BUFX2 g_N3343 (N626, N3343);
	AND2X1 g_N3344 (N1347, N567, N3344);
	INVX1 g_N3345 (N2951, N3345);
	BUFX2 g_N357 (N2653, N357);
	BUFX2 g_N3346 (N2362, N3346);
	INVX1 g_N3347 (N3828, N3347);
	BUFX2 g_N3348 (N892, N3348);
	BUFX2 g_N3349 (N1037, N3349);
	BUFX2 g_N3350 (N2593, N3350);
	INVX1 g_N3351 (N1112, N3351);
	AND2X1 g_N3352 (N3176, N2687, N3352);
	BUFX2 g_N3353 (N2722, N3353);
	INVX1 g_N3354 (N1119, N3354);
	BUFX2 g_N3355 (N3127, N3355);
	BUFX2 g_N3356 (N3799, N3356);
	INVX1 g_N3357 (N1085, N3357);
	INVX1 g_N3358 (N2877, N3358);
	INVX1 g_N3359 (N32, N3359);
	AND2X1 g_N3360 (N3452, N1628, N3360);
	BUFX2 g_N3361 (N1462, N3361);
	INVX1 g_N3362 (N2387, N3362);
	INVX1 g_N3363 (N2315, N3363);
	BUFX2 g_N3364 (N3557, N3364);
	BUFX2 g_N3365 (N603, N3365);
	AND2X1 g_N3366 (N3758, N823, N3366);
	BUFX2 g_N3367 (N2797, N3367);
	BUFX2 g_N3368 (N2789, N3368);
	INVX1 g_N3369 (N3330, N3369);
	INVX1 g_N3370 (N3739, N3370);
	BUFX2 g_N3371 (N3695, N3371);
	AND2X1 g_N3372 (N2654, N3818, N3372);
	INVX1 g_N3373 (N2870, N3373);
	INVX1 g_N3374 (N1468, N3374);
	AND2X1 g_N3375 (N1418, N1896, N3375);
	BUFX2 g_N3376 (N3186, N3376);
	BUFX2 g_N3377 (N3500, N3377);
	INVX1 g_N3378 (N1200, N3378);
	INVX1 g_N3379 (N2733, N3379);
	AND2X1 g_N3380 (N2283, N2469, N3380);
	INVX1 g_N3381 (N1682, N3381);
	AND2X1 g_N3382 (N1078, N2829, N3382);
	AND2X1 g_N3383 (N2723, N1377, N3383);
	INVX1 g_N3384 (N2656, N3384);
	BUFX2 g_N3385 (N3230, N3385);
	BUFX2 g_N3386 (N2343, N3386);
	INVX1 g_N3387 (N1550, N3387);
	INVX1 g_N3388 (N2798, N3388);
	BUFX2 g_N3389 (N1053, N3389);
	AND2X1 g_N3390 (N66, N119, N3390);
	BUFX2 g_N3391 (N3829, N3391);
	AND2X1 g_N3392 (N2832, N3794, N3392);
	BUFX2 g_N3393 (N898, N3393);
	INVX1 g_N3394 (N1517, N3394);
	BUFX2 g_N3395 (N1631, N3395);
	BUFX2 g_N3396 (N1593, N3396);
	INVX1 g_N3397 (N3335, N3397);
	AND2X1 g_N3398 (N3042, N2258, N3398);
	INVX1 g_N3399 (N3674, N3399);
	INVX1 g_N3400 (N3059, N3400);
	BUFX2 g_N358 (N2514, N358);
	AND2X1 g_N3401 (N1137, N3499, N3401);
	BUFX2 g_N3402 (N2308, N3402);
	BUFX2 g_N3403 (N3261, N3403);
	INVX1 g_N3404 (N2894, N3404);
	AND2X1 g_N3405 (N2957, N2596, N3405);
	INVX1 g_N3406 (N127, N3406);
	BUFX2 g_N3407 (N3089, N3407);
	AND2X1 g_N3408 (N2741, N2072, N3408);
	BUFX2 g_N3409 (N2658, N3409);
	BUFX2 g_N3410 (N3443, N3410);
	INVX1 g_N3411 (N781, N3411);
	AND2X1 g_N3412 (N431, N3011, N3412);
	INVX1 g_N3413 (N1697, N3413);
	AND2X1 g_N3414 (N2567, N605, N3414);
	INVX1 g_N3415 (N2144, N3415);
	AND2X1 g_N3416 (N393, N3470, N3416);
	AND2X1 g_N3417 (N2432, N3378, N3417);
	INVX1 g_N3418 (N1259, N3418);
	BUFX2 g_N3419 (N1888, N3419);
	BUFX2 g_N3420 (N3522, N3420);
	INVX1 g_N3421 (N2861, N3421);
	BUFX2 g_N3422 (N1475, N3422);
	AND2X1 g_N3423 (N2297, N1556, N3423);
	INVX1 g_N3424 (N1146, N3424);
	INVX1 g_N3425 (N3588, N3425);
	INVX1 g_N3426 (N879, N3426);
	INVX1 g_N3427 (N1293, N3427);
	BUFX2 g_N3428 (N2365, N3428);
	AND2X1 g_N3429 (N3291, N3920, N3429);
	INVX1 g_N3430 (N1964, N3430);
	INVX1 g_N3431 (N20, N3431);
	BUFX2 g_N3432 (N412, N3432);
	BUFX2 g_N3433 (N2095, N3433);
	BUFX2 g_N3434 (N2745, N3434);
	AND2X1 g_N3435 (N407, N2349, N3435);
	BUFX2 g_N3436 (N3830, N3436);
	BUFX2 g_N3437 (N1401, N3437);
	INVX1 g_N3438 (N2430, N3438);
	INVX1 g_N3439 (N3891, N3439);
	INVX1 g_N3440 (N3117, N3440);
	INVX1 g_N3441 (N240, N3441);
	BUFX2 g_N359 (N2563, N359);
	INVX1 g_N3442 (N2860, N3442);
	AND2X1 g_N3443 (N1492, N3653, N3443);
	AND2X1 g_N3444 (N3782, N2085, N3444);
	AND2X1 g_N3445 (N3233, N468, N3445);
	AND2X1 g_N3446 (N3870, N2458, N3446);
	BUFX2 g_N360 (N3395, N360);
	BUFX2 g_N3447 (N3197, N3447);
	AND2X1 g_N3448 (N3697, N3413, N3448);
	BUFX2 g_N3449 (N2476, N3449);
	BUFX2 g_N3450 (N1519, N3450);
	BUFX2 g_N361 (N2605, N361);
	INVX1 g_N3451 (N2142, N3451);
	BUFX2 g_N362 (N522, N362);
	INVX1 g_N3452 (N2152, N3452);
	BUFX2 g_N3453 (N3405, N3453);
	INVX1 g_N3454 (N7, N3454);
	AND2X1 g_N3455 (N2779, N3234, N3455);
	AND2X1 g_N3456 (N1148, N3643, N3456);
	INVX1 g_N3457 (N1314, N3457);
	INVX1 g_N3458 (N2948, N3458);
	AND2X1 g_N3459 (N165, N31, N3459);
	AND2X1 g_N3460 (N150, N101, N3460);
	AND2X1 g_N3461 (N1090, N627, N3461);
	AND2X1 g_N3462 (N3481, N989, N3462);
	BUFX2 g_N3463 (N1360, N3463);
	BUFX2 g_N3464 (N2457, N3464);
	INVX1 g_N3465 (N2306, N3465);
	BUFX2 g_N3466 (N1952, N3466);
	AND2X1 g_N3467 (N3667, N1233, N3467);
	BUFX2 g_N363 (N3349, N363);
	AND2X1 g_N3468 (N1815, N3792, N3468);
	INVX1 g_N3469 (N3503, N3469);
	BUFX2 g_N3470 (N3073, N3470);
	AND2X1 g_N3471 (N3548, N3098, N3471);
	INVX1 g_N3472 (N615, N3472);
	AND2X1 g_N3473 (N3668, N2120, N3473);
	INVX1 g_N3474 (N622, N3474);
	AND2X1 g_N3475 (N631, N2742, N3475);
	INVX1 g_N3476 (N2931, N3476);
	INVX1 g_N3477 (N3322, N3477);
	BUFX2 g_N3478 (N1036, N3478);
	INVX1 g_N3479 (N78, N3479);
	AND2X1 g_N3480 (N3560, N3241, N3480);
	INVX1 g_N3481 (N3749, N3481);
	AND2X1 g_N3482 (N1574, N2984, N3482);
	INVX1 g_N3483 (N2165, N3483);
	INVX1 g_N3484 (N1077, N3484);
	INVX1 g_N3485 (N997, N3485);
	INVX1 g_N3486 (N2645, N3486);
	AND2X1 g_N3487 (N2522, N541, N3487);
	BUFX2 g_N3488 (N630, N3488);
	BUFX2 g_N3489 (N3398, N3489);
	AND2X1 g_N3490 (N2461, N3669, N3490);
	BUFX2 g_N3491 (N2665, N3491);
	BUFX2 g_N3492 (N3874, N3492);
	AND2X1 g_N3493 (N3788, N1265, N3493);
	AND2X1 g_N3494 (N3164, N1741, N3494);
	INVX1 g_N3495 (N2744, N3495);
	INVX1 g_N3496 (N3850, N3496);
	INVX1 g_N3497 (N2262, N3497);
	AND2X1 g_N3498 (N2225, N2692, N3498);
	INVX1 g_N3499 (N3149, N3499);
	AND2X1 g_N3500 (N3379, N3937, N3500);
	INVX1 g_N3501 (N443, N3501);
	BUFX2 g_N3502 (N3708, N3502);
	BUFX2 g_N3503 (N2987, N3503);
	BUFX2 g_N3504 (N1907, N3504);
	BUFX2 g_N3505 (N1799, N3505);
	AND2X1 g_N3506 (N3875, N2799, N3506);
	INVX1 g_N3507 (N137, N3507);
	INVX1 g_N3508 (N580, N3508);
	INVX1 g_N3509 (N1317, N3509);
	INVX1 g_N3510 (N3899, N3510);
	BUFX2 g_N3511 (N1061, N3511);
	INVX1 g_N3512 (N2203, N3512);
	INVX1 g_N3513 (N46, N3513);
	AND2X1 g_N3514 (N782, N753, N3514);
	BUFX2 g_N3515 (N2521, N3515);
	AND2X1 g_N3516 (N1634, N2846, N3516);
	AND2X1 g_N3517 (N218, N33, N3517);
	INVX1 g_N3518 (N87, N3518);
	BUFX2 g_N364 (N639, N364);
	INVX1 g_N3519 (N3269, N3519);
	INVX1 g_N3520 (N2325, N3520);
	AND2X1 g_N3521 (N3458, N3725, N3521);
	AND2X1 g_N3522 (N1504, N3001, N3522);
	AND2X1 g_N3523 (N795, N1779, N3523);
	BUFX2 g_N3524 (N1339, N3524);
	AND2X1 g_N3525 (N1531, N3250, N3525);
	AND2X1 g_N3526 (N1782, N871, N3526);
	AND2X1 g_N3527 (N2108, N767, N3527);
	BUFX2 g_N365 (N2855, N365);
	BUFX2 g_N3528 (N3521, N3528);
	INVX1 g_N3529 (N2547, N3529);
	AND2X1 g_N3530 (N3107, N766, N3530);
	BUFX2 g_N3531 (N3832, N3531);
	BUFX2 g_N3532 (N1686, N3532);
	AND2X1 g_N3533 (N3064, N2218, N3533);
	AND2X1 g_N3534 (N2026, N2094, N3534);
	BUFX2 g_N3535 (N851, N3535);
	BUFX2 g_N3536 (N1724, N3536);
	INVX1 g_N3537 (N524, N3537);
	BUFX2 g_N366 (N3063, N366);
	AND2X1 g_N3538 (N3472, N2673, N3538);
	AND2X1 g_N3539 (N2794, N2628, N3539);
	BUFX2 g_N3540 (N1214, N3540);
	BUFX2 g_N3541 (N2081, N3541);
	BUFX2 g_N367 (N1871, N367);
	INVX1 g_N3542 (N3450, N3542);
	BUFX2 g_N3543 (N807, N3543);
	INVX1 g_N3544 (N2550, N3544);
	BUFX2 g_N3545 (N3459, N3545);
	INVX1 g_N3546 (N3504, N3546);
	AND2X1 g_N3547 (N2230, N2383, N3547);
	BUFX2 g_N3548 (N2824, N3548);
	BUFX2 g_N3549 (N641, N3549);
	INVX1 g_N3550 (N1842, N3550);
	AND2X1 g_N3551 (N2889, N446, N3551);
	INVX1 g_N3552 (N2646, N3552);
	INVX1 g_N3553 (N2614, N3553);
	INVX1 g_N3554 (N1830, N3554);
	INVX1 g_N3555 (N3819, N3555);
	BUFX2 g_N3556 (N3493, N3556);
	AND2X1 g_N3557 (N2639, N1091, N3557);
	BUFX2 g_N3558 (N3898, N3558);
	BUFX2 g_N3559 (N1123, N3559);
	INVX1 g_N3560 (N2259, N3560);
	BUFX2 g_N3561 (N3244, N3561);
	INVX1 g_N3562 (N1235, N3562);
	INVX1 g_N3563 (N2134, N3563);
	BUFX2 g_N3564 (N1664, N3564);
	AND2X1 g_N3565 (N950, N495, N3565);
	INVX1 g_N3566 (N1181, N3566);
	AND2X1 g_N3567 (N118, N158, N3567);
	AND2X1 g_N3568 (N3705, N2953, N3568);
	AND2X1 g_N3569 (N2281, N3044, N3569);
	INVX1 g_N3570 (N219, N3570);
	INVX1 g_N3571 (N41, N3571);
	AND2X1 g_N3572 (N2691, N492, N3572);
	BUFX2 g_N3573 (N1118, N3573);
	AND2X1 g_N3574 (N2633, N1805, N3574);
	BUFX2 g_N3575 (N1143, N3575);
	BUFX2 g_N3576 (N737, N3576);
	INVX1 g_N3577 (N2952, N3577);
	AND2X1 g_N3578 (N913, N1849, N3578);
	INVX1 g_N3579 (N52, N3579);
	BUFX2 g_N3580 (N2657, N3580);
	INVX1 g_N3581 (N2518, N3581);
	INVX1 g_N3582 (N778, N3582);
	BUFX2 g_N3583 (N3372, N3583);
	INVX1 g_N3584 (N2560, N3584);
	INVX1 g_N3585 (N2241, N3585);
	INVX1 g_N3586 (N1770, N3586);
	INVX1 g_N3587 (N3749, N3587);
	BUFX2 g_N3588 (N2881, N3588);
	INVX1 g_N3589 (N3556, N3589);
	INVX1 g_N3590 (N1258, N3590);
	BUFX2 g_N3591 (N1978, N3591);
	INVX1 g_N3592 (N1407, N3592);
	BUFX2 g_N3593 (N3894, N3593);
	BUFX2 g_N3594 (N3498, N3594);
	BUFX2 g_N3595 (N2876, N3595);
	INVX1 g_N3596 (N889, N3596);
	INVX1 g_N3597 (N180, N3597);
	INVX1 g_N3598 (N1487, N3598);
	INVX1 g_N3599 (N174, N3599);
	INVX1 g_N3600 (N392, N3600);
	INVX1 g_N3601 (N2024, N3601);
	AND2X1 g_N3602 (N3621, N1858, N3602);
	INVX1 g_N3603 (N170, N3603);
	INVX1 g_N3604 (N454, N3604);
	AND2X1 g_N3605 (N240, N50, N3605);
	INVX1 g_N3606 (N3807, N3606);
	INVX1 g_N3607 (N1003, N3607);
	AND2X1 g_N3608 (N2199, N2028, N3608);
	INVX1 g_N3609 (N1176, N3609);
	INVX1 g_N3610 (N2411, N3610);
	AND2X1 g_N3611 (N1571, N3108, N3611);
	INVX1 g_N3612 (N1322, N3612);
	BUFX2 g_N368 (N3071, N368);
	BUFX2 g_N3613 (N3423, N3613);
	BUFX2 g_N3614 (N3101, N3614);
	BUFX2 g_N3615 (N1506, N3615);
	INVX1 g_N3616 (N1228, N3616);
	INVX1 g_N3617 (N29, N3617);
	AND2X1 g_N3618 (N1966, N1909, N3618);
	BUFX2 g_N3619 (N2139, N3619);
	INVX1 g_N3620 (N2807, N3620);
	INVX1 g_N3621 (N713, N3621);
	INVX1 g_N3622 (N209, N3622);
	AND2X1 g_N3623 (N3327, N735, N3623);
	AND2X1 g_N3624 (N254, N207, N3624);
	BUFX2 g_N369 (N1313, N369);
	INVX1 g_N3625 (N164, N3625);
	INVX1 g_N3626 (N1354, N3626);
	BUFX2 g_N3627 (N1719, N3627);
	BUFX2 g_N3628 (N2878, N3628);
	BUFX2 g_N3629 (N3446, N3629);
	INVX1 g_N3630 (N3545, N3630);
	BUFX2 g_N3631 (N3578, N3631);
	INVX1 g_N3632 (N1170, N3632);
	INVX1 g_N3633 (N44, N3633);
	BUFX2 g_N3634 (N3897, N3634);
	BUFX2 g_N3635 (N1737, N3635);
	BUFX2 g_N3636 (N2351, N3636);
	AND2X1 g_N3637 (N197, N88, N3637);
	INVX1 g_N3638 (N136, N3638);
	INVX1 g_N3639 (N84, N3639);
	INVX1 g_N3640 (N24, N3640);
	BUFX2 g_N3641 (N2016, N3641);
	AND2X1 g_N3642 (N1298, N2397, N3642);
	INVX1 g_N3643 (N2224, N3643);
	INVX1 g_N3644 (N3593, N3644);
	BUFX2 g_N3645 (N1386, N3645);
	INVX1 g_N3646 (N1592, N3646);
	BUFX2 g_N370 (N1524, N370);
	BUFX2 g_N3647 (N588, N3647);
	INVX1 g_N3648 (N1684, N3648);
	BUFX2 g_N3649 (N3795, N3649);
	INVX1 g_N3650 (N1046, N3650);
	INVX1 g_N3651 (N3117, N3651);
	INVX1 g_N3652 (N1867, N3652);
	INVX1 g_N3653 (N1440, N3653);
	BUFX2 g_N3654 (N1833, N3654);
	AND2X1 g_N3655 (N2697, N949, N3655);
	BUFX2 g_N3656 (N3161, N3656);
	INVX1 g_N3657 (N2377, N3657);
	INVX1 g_N3658 (N1729, N3658);
	INVX1 g_N3659 (N1413, N3659);
	INVX1 g_N3660 (N1674, N3660);
	AND2X1 g_N3661 (N107, N103, N3661);
	AND2X1 g_N3662 (N1876, N3909, N3662);
	BUFX2 g_N3663 (N2321, N3663);
	INVX1 g_N3664 (N997, N3664);
	AND2X1 g_N3665 (N3801, N1505, N3665);
	INVX1 g_N3666 (N59, N3666);
	INVX1 g_N3667 (N2995, N3667);
	BUFX2 g_N3668 (N3490, N3668);
	INVX1 g_N3669 (N3559, N3669);
	INVX1 g_N3670 (N3777, N3670);
	AND2X1 g_N3671 (N1282, N2465, N3671);
	BUFX2 g_N3672 (N2703, N3672);
	BUFX2 g_N3673 (N729, N3673);
	BUFX2 g_N3674 (N1311, N3674);
	AND2X1 g_N3675 (N3054, N1915, N3675);
	INVX1 g_N3676 (N3466, N3676);
	INVX1 g_N3677 (N3277, N3677);
	INVX1 g_N3678 (N1219, N3678);
	AND2X1 g_N3679 (N1637, N2726, N3679);
	INVX1 g_N3680 (N1535, N3680);
	INVX1 g_N3681 (N2747, N3681);
	INVX1 g_N3682 (N182, N3682);
	AND2X1 g_N3683 (N3585, N916, N3683);
	BUFX2 g_N3684 (N1182, N3684);
	BUFX2 g_N3685 (N1918, N3685);
	INVX1 g_N3686 (N1022, N3686);
	INVX1 g_N3687 (N1899, N3687);
	INVX1 g_N3688 (N2838, N3688);
	INVX1 g_N3689 (N95, N3689);
	AND2X1 g_N3690 (N43, N64, N3690);
	INVX1 g_N3691 (N2609, N3691);
	BUFX2 g_N371 (N2752, N371);
	INVX1 g_N3692 (N3515, N3692);
	INVX1 g_N3693 (N3312, N3693);
	INVX1 g_N3694 (N675, N3694);
	AND2X1 g_N3695 (N2569, N3333, N3695);
	INVX1 g_N3696 (N1603, N3696);
	INVX1 g_N3697 (N1681, N3697);
	AND2X1 g_N3698 (N3687, N3691, N3698);
	BUFX2 g_N3699 (N3344, N3699);
	BUFX2 g_N3700 (N1324, N3700);
	BUFX2 g_N372 (N570, N372);
	AND2X1 g_N3701 (N1689, N387, N3701);
	OR2X1 g_N3702 (N3636, N3396, N3702);
	AND2X1 g_N3703 (N3166, N781, N3703);
	AND2X1 g_N3704 (N3424, N1052, N3704);
	INVX1 g_N3705 (N408, N3705);
	AND2X1 g_N3706 (N1336, N2334, N3706);
	AND2X1 g_N3707 (N2976, N2174, N3707);
	AND2X1 g_N3708 (N26, N252, N3708);
	AND2X1 g_N3709 (N3660, N2441, N3709);
	BUFX2 g_N3710 (N3750, N3710);
	INVX1 g_N3711 (N3685, N3711);
	BUFX2 g_N373 (N1291, N373);
	BUFX2 g_N3712 (N2866, N3712);
	BUFX2 g_N3713 (N979, N3713);
	BUFX2 g_N3714 (N1941, N3714);
	BUFX2 g_N3715 (N1804, N3715);
	INVX1 g_N3716 (N3536, N3716);
	BUFX2 g_N3717 (N594, N3717);
	AND2X1 g_N3718 (N3563, N2597, N3718);
	INVX1 g_N3719 (N3714, N3719);
	AND2X1 g_N3720 (N3699, N1202, N3720);
	BUFX2 g_N3721 (N728, N3721);
	AND2X1 g_N3722 (N2330, N2972, N3722);
	BUFX2 g_N3723 (N2882, N3723);
	BUFX2 g_N374 (N3391, N374);
	INVX1 g_N3724 (N1119, N3724);
	BUFX2 g_N375 (N2435, N375);
	INVX1 g_N3725 (N904, N3725);
	AND2X1 g_N3726 (N1863, N1207, N3726);
	AND2X1 g_N3727 (N1927, N1180, N3727);
	BUFX2 g_N3728 (N2237, N3728);
	INVX1 g_N3729 (N2542, N3729);
	INVX1 g_N3730 (N2105, N3730);
	INVX1 g_N3731 (N520, N3731);
	INVX1 g_N3732 (N1527, N3732);
	INVX1 g_N3733 (N2286, N3733);
	INVX1 g_N3734 (N2922, N3734);
	INVX1 g_N3735 (N125, N3735);
	INVX1 g_N3736 (N1751, N3736);
	INVX1 g_N3737 (N3940, N3737);
	BUFX2 g_N3738 (N3016, N3738);
	BUFX2 g_N3739 (N2221, N3739);
	INVX1 g_N3740 (N205, N3740);
	AND2X1 g_N3741 (N2352, N2302, N3741);
	INVX1 g_N3742 (N94, N3742);
	INVX1 g_N3743 (N3409, N3743);
	AND2X1 g_N3744 (N3404, N3652, N3744);
	BUFX2 g_N3745 (N1714, N3745);
	BUFX2 g_N3746 (N2301, N3746);
	INVX1 g_N3747 (N443, N3747);
	INVX1 g_N3748 (N118, N3748);
	BUFX2 g_N3749 (N2223, N3749);
	AND2X1 g_N3750 (N2194, N2676, N3750);
	BUFX2 g_N3751 (N3221, N3751);
	INVX1 g_N3752 (N1402, N3752);
	INVX1 g_N3753 (N582, N3753);
	AND2X1 g_N3754 (N3265, N684, N3754);
	AND2X1 g_N3755 (N2989, N1660, N3755);
	BUFX2 g_N376 (N2217, N376);
	INVX1 g_N3756 (N2240, N3756);
	AND2X1 g_N3757 (N2235, N1390, N3757);
	INVX1 g_N3758 (N391, N3758);
	AND2X1 g_N3759 (N2141, N3397, N3759);
	AND2X1 g_N3760 (N138, N212, N3760);
	INVX1 g_N3761 (N3805, N3761);
	INVX1 g_N3762 (N1340, N3762);
	AND2X1 g_N3763 (N3537, N2305, N3763);
	BUFX2 g_N3764 (N863, N3764);
	AND2X1 g_N3765 (N2445, N1327, N3765);
	BUFX2 g_N377 (N1777, N377);
	AND2X1 g_N3766 (N3743, N2659, N3766);
	BUFX2 g_N3767 (N794, N3767);
	AND2X1 g_N3768 (N1050, N2419, N3768);
	AND2X1 g_N3769 (N3433, N2303, N3769);
	INVX1 g_N3770 (N1902, N3770);
	INVX1 g_N3771 (N2702, N3771);
	INVX1 g_N3772 (N3854, N3772);
	AND2X1 g_N3773 (N1114, N2339, N3773);
	INVX1 g_N3774 (N2640, N3774);
	INVX1 g_N3775 (N3715, N3775);
	AND2X1 g_N3776 (N1879, N2729, N3776);
	BUFX2 g_N3777 (N2453, N3777);
	INVX1 g_N3778 (N1272, N3778);
	BUFX2 g_N3779 (N822, N3779);
	INVX1 g_N3780 (N3327, N3780);
	AND2X1 g_N3781 (N1850, N1621, N3781);
	BUFX2 g_N3782 (N2787, N3782);
	INVX1 g_N3783 (N2418, N3783);
	INVX1 g_N3784 (N89, N3784);
	AND2X1 g_N3785 (N1394, N997, N3785);
	INVX1 g_N3786 (N2581, N3786);
	INVX1 g_N3787 (N554, N3787);
	INVX1 g_N3788 (N3877, N3788);
	INVX1 g_N3789 (N69, N3789);
	AND2X1 g_N3790 (N2119, N1405, N3790);
	BUFX2 g_N3791 (N860, N3791);
	INVX1 g_N3792 (N2369, N3792);
	BUFX2 g_N3793 (N867, N3793);
	INVX1 g_N3794 (N121, N3794);
	AND2X1 g_N3795 (N1367, N3780, N3795);
	AND2X1 g_N3796 (N255, N72, N3796);
	INVX1 g_N3797 (N1802, N3797);
	INVX1 g_N3798 (N3018, N3798);
	AND2X1 g_N3799 (N3266, N1555, N3799);
	BUFX2 g_N3800 (N803, N3800);
	INVX1 g_N3801 (N910, N3801);
	BUFX2 g_N3802 (N1608, N3802);
	INVX1 g_N3803 (N2388, N3803);
	AND2X1 g_N3804 (N123, N191, N3804);
	BUFX2 g_N3805 (N1652, N3805);
	AND2X1 g_N3806 (N3278, N685, N3806);
	BUFX2 g_N3807 (N2604, N3807);
	INVX1 g_N3808 (N1430, N3808);
	AND2X1 g_N3809 (N1126, N459, N3809);
	INVX1 g_N3810 (N1647, N3810);
	INVX1 g_N3811 (N2623, N3811);
	BUFX2 g_N3812 (N577, N3812);
	AND2X1 g_N3813 (N3105, N1642, N3813);
	INVX1 g_N3814 (N1375, N3814);
	INVX1 g_N3815 (N1628, N3815);
	BUFX2 g_N3816 (N1818, N3816);
	AND2X1 g_N3817 (N2214, N2535, N3817);
	INVX1 g_N3818 (N1925, N3818);
	BUFX2 g_N3819 (N1735, N3819);
	AND2X1 g_N3820 (N3354, N3357, N3820);
	BUFX2 g_N3821 (N2442, N3821);
	AND2X1 g_N3822 (N1544, N3552, N3822);
	BUFX2 g_N378 (N1522, N378);
	INVX1 g_N3823 (N63, N3823);
	INVX1 g_N3824 (N3575, N3824);
	AND2X1 g_N3825 (N3910, N1385, N3825);
	AND2X1 g_N3826 (N3753, N576, N3826);
	INVX1 g_N3827 (N1112, N3827);
	BUFX2 g_N3828 (N3444, N3828);
	AND2X1 g_N3829 (N696, N2991, N3829);
	AND2X1 g_N3830 (N2776, N3053, N3830);
	INVX1 g_N3831 (N2411, N3831);
	AND2X1 g_N3832 (N2526, N2097, N3832);
	INVX1 g_N3833 (N2314, N3833);
	BUFX2 g_N3834 (N3471, N3834);
	AND2X1 g_N3835 (N1806, N3008, N3835);
	BUFX2 g_N3836 (N2003, N3836);
	BUFX2 g_N3837 (N948, N3837);
	BUFX2 g_N3838 (N1201, N3838);
	INVX1 g_N3839 (N2503, N3839);
	BUFX2 g_N379 (N1832, N379);
	BUFX2 g_N3840 (N1635, N3840);
	BUFX2 g_N3841 (N742, N3841);
	INVX1 g_N3842 (N2509, N3842);
	AND2X1 g_N3843 (N2879, N421, N3843);
	INVX1 g_N3844 (N3909, N3844);
	AND2X1 g_N3845 (N669, N1286, N3845);
	BUFX2 g_N380 (N2008, N380);
	INVX1 g_N3846 (N64, N3846);
	AND2X1 g_N3847 (N3104, N968, N3847);
	INVX1 g_N3848 (N2, N3848);
	AND2X1 g_N3849 (N1345, N3562, N3849);
	BUFX2 g_N3850 (N883, N3850);
	INVX1 g_N3851 (N2737, N3851);
	AND2X1 g_N3852 (N1890, N3504, N3852);
	INVX1 g_N3853 (N3293, N3853);
	BUFX2 g_N3854 (N3776, N3854);
	INVX1 g_N3855 (N518, N3855);
	AND2X1 g_N3856 (N3586, N706, N3856);
	INVX1 g_N3857 (N228, N3857);
	BUFX2 g_N3858 (N3338, N3858);
	INVX1 g_N3859 (N39, N3859);
	AND2X1 g_N3860 (N69, N19, N3860);
	INVX1 g_N3861 (N2158, N3861);
	INVX1 g_N3862 (N2420, N3862);
	INVX1 g_N3863 (N2500, N3863);
	BUFX2 g_N3864 (N2460, N3864);
	AND2X1 g_N3865 (N978, N1258, N3865);
	INVX1 g_N3866 (N2951, N3866);
	BUFX2 g_N3867 (N727, N3867);
	INVX1 g_N3868 (N233, N3868);
	AND2X1 g_N3869 (N1262, N2805, N3869);
	INVX1 g_N3870 (N2196, N3870);
	BUFX2 g_N3871 (N1680, N3871);
	INVX1 g_N3872 (N483, N3872);
	AND2X1 g_N3873 (N3544, N1729, N3873);
	AND2X1 g_N3874 (N2929, N3271, N3874);
	INVX1 g_N3875 (N747, N3875);
	INVX1 g_N3876 (N93, N3876);
	BUFX2 g_N3877 (N3523, N3877);
	INVX1 g_N3878 (N148, N3878);
	AND2X1 g_N3879 (N1541, N700, N3879);
	INVX1 g_N3880 (N248, N3880);
	AND2X1 g_N3881 (N56, N156, N3881);
	BUFX2 g_N3882 (N1648, N3882);
	AND2X1 g_N3883 (N1919, N1693, N3883);
	BUFX2 g_N3884 (N817, N3884);
	BUFX2 g_N381 (N2327, N381);
	INVX1 g_N3885 (N2057, N3885);
	BUFX2 g_N3886 (N2710, N3886);
	BUFX2 g_N3887 (N1655, N3887);
	BUFX2 g_N3888 (N610, N3888);
	INVX1 g_N3889 (N3156, N3889);
	AND2X1 g_N3890 (N55, N29, N3890);
	BUFX2 g_N3891 (N3417, N3891);
	BUFX2 g_N3892 (N2828, N3892);
	INVX1 g_N3893 (N2836, N3893);
	BUFX2 g_N382 (N1986, N382);
	AND2X1 g_N3894 (N2777, N2920, N3894);
	INVX1 g_N3895 (N2384, N3895);
	INVX1 g_N3896 (N2920, N3896);
	AND2X1 g_N3897 (N1318, N1017, N3897);
	AND2X1 g_N3898 (N1330, N3606, N3898);
	BUFX2 g_N3899 (N2539, N3899);
	BUFX2 g_N3900 (N606, N3900);
	AND2X1 g_N3901 (N2378, N3259, N3901);
	BUFX2 g_N3902 (N1369, N3902);
	BUFX2 g_N3903 (N2763, N3903);
	AND2X1 g_N3904 (N590, N2758, N3904);
	INVX1 g_N3905 (N3314, N3905);
	BUFX2 g_N3906 (N3321, N3906);
	AND2X1 g_N3907 (N549, N3577, N3907);
	INVX1 g_N3908 (N595, N3908);
	BUFX2 g_N3909 (N3475, N3909);
	INVX1 g_N3910 (N654, N3910);
	AND2X1 g_N3911 (N2272, N2036, N3911);
	BUFX2 g_N3912 (N1393, N3912);
	INVX1 g_N3913 (N3887, N3913);
	AND2X1 g_N3914 (N1982, N1512, N3914);
	BUFX2 g_N3915 (N514, N3915);
	BUFX2 g_N3916 (N3611, N3916);
	INVX1 g_N3917 (N1800, N3917);
	BUFX2 g_N3918 (N811, N3918);
	AND2X1 g_N3919 (N231, N251, N3919);
	INVX1 g_N3920 (N1328, N3920);
	AND2X1 g_N3921 (N1883, N2440, N3921);
	INVX1 g_N3922 (N17, N3922);
	AND2X1 g_N3923 (N723, N3601, N3923);
	INVX1 g_N3924 (N3036, N3924);
	AND2X1 g_N3925 (N59, N168, N3925);
	INVX1 g_N3926 (N2434, N3926);
	BUFX2 g_N3927 (N2073, N3927);
	AND2X1 g_N3928 (N144, N185, N3928);
	AND2X1 g_N3929 (N2079, N1763, N3929);
	AND2X1 g_N3930 (N3255, N620, N3930);
	BUFX2 g_N3931 (N1373, N3931);
	INVX1 g_N3932 (N2599, N3932);
	BUFX2 g_N3933 (N2192, N3933);
	INVX1 g_N3934 (N1765, N3934);
	INVX1 g_N3935 (N1983, N3935);
	AND2X1 g_N3936 (N3737, N531, N3936);
	BUFX2 g_N383 (N3812, N383);
	INVX1 g_N3937 (N3055, N3937);
	BUFX2 g_N3938 (N3065, N3938);
	BUFX2 g_N3939 (N3928, N3939);
	BUFX2 g_N3940 (N2667, N3940);
	INVX1 g_N3941 (N3464, N3941);
	INVX1 g_N3942 (N3292, N3942);
	AND2X1 g_N3943 (N3733, N2088, N3943);
	BUFX2 g_N384 (N3279, N384);
	BUFX2 g_N385 (N2410, N385);
	INVX1 g_N3944 (N3654, N3944);
	INVX1 g_N3945 (N2809, N3945);
	BUFX2 g_N3946 (N2228, N3946);

endmodule
